library verilog;
use verilog.vl_types.all;
entity FIR_avr_tst is
end FIR_avr_tst;
