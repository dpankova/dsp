////////////////////////////////////////////////////////////////
// Daria Pankova Wed Jul 22 12:20:07 EDT 2015
// test_rom.v
//
// "Pseudo RAM with baseline data"
// A custom Verilog HDL module.
// 
////////////////////////////////////////////////////////////////


module test_rom_example(
		input [12:0]   rdaddr,
		output [13:0] adc_val
		);
   reg [13:0] adc_rom[0:6778];
   
   assign adc_val = adc_rom[rdaddr];
   
   initial begin
      adc_rom[0] <= 8185;
      adc_rom[1] <= 8185;
      adc_rom[2] <= 8187;
      adc_rom[3] <= 8187;
      adc_rom[4] <= 8186;
      adc_rom[5] <= 8185;
      adc_rom[6] <= 8187;
      adc_rom[7] <= 8185;
      adc_rom[8] <= 8187;
      adc_rom[9] <= 8186;
      adc_rom[10] <= 8185;
      adc_rom[11] <= 8186;
      adc_rom[12] <= 8187;
      adc_rom[13] <= 8184;
      adc_rom[14] <= 8186;
      adc_rom[15] <= 8186;
      adc_rom[16] <= 8185;
      adc_rom[17] <= 8186;
      adc_rom[18] <= 8186;
      adc_rom[19] <= 8187;
      adc_rom[20] <= 8186;
      adc_rom[21] <= 8185;
      adc_rom[22] <= 8185;
      adc_rom[23] <= 8183;
      adc_rom[24] <= 8187;
      adc_rom[25] <= 8183;
      adc_rom[26] <= 8186;
      adc_rom[27] <= 8187;
      adc_rom[28] <= 8185;
      adc_rom[29] <= 8187;
      adc_rom[30] <= 8186;
      adc_rom[31] <= 8187;
      adc_rom[32] <= 8185;
      adc_rom[33] <= 8184;
      adc_rom[34] <= 8187;
      adc_rom[35] <= 8187;
      adc_rom[36] <= 8185;
      adc_rom[37] <= 8187;
      adc_rom[38] <= 8185;
      adc_rom[39] <= 8188;
      adc_rom[40] <= 8187;
      adc_rom[41] <= 8186;
      adc_rom[42] <= 8189;
      adc_rom[43] <= 8186;
      adc_rom[44] <= 8188;
      adc_rom[45] <= 8185;
      adc_rom[46] <= 8186;
      adc_rom[47] <= 8188;
      adc_rom[48] <= 8186;
      adc_rom[49] <= 8186;
      adc_rom[50] <= 8186;
      adc_rom[51] <= 8187;
      adc_rom[52] <= 8186;
      adc_rom[53] <= 8185;
      adc_rom[54] <= 8187;
      adc_rom[55] <= 8185;
      adc_rom[56] <= 8186;
      adc_rom[57] <= 8187;
      adc_rom[58] <= 8187;
      adc_rom[59] <= 8186;
      adc_rom[60] <= 8186;
      adc_rom[61] <= 8186;
      adc_rom[62] <= 8188;
      adc_rom[63] <= 8186;
      adc_rom[64] <= 8186;
      adc_rom[65] <= 8186;
      adc_rom[66] <= 8188;
      adc_rom[67] <= 8186;
      adc_rom[68] <= 8185;
      adc_rom[69] <= 8188;
      adc_rom[70] <= 8186;
      adc_rom[71] <= 8188;
      adc_rom[72] <= 8187;
      adc_rom[73] <= 8185;
      adc_rom[74] <= 8188;
      adc_rom[75] <= 8187;
      adc_rom[76] <= 8186;
      adc_rom[77] <= 8188;
      adc_rom[78] <= 8184;
      adc_rom[79] <= 8189;
      adc_rom[80] <= 8187;
      adc_rom[81] <= 8186;
      adc_rom[82] <= 8185;
      adc_rom[83] <= 8183;
      adc_rom[84] <= 8189;
      adc_rom[85] <= 8185;
      adc_rom[86] <= 8188;
      adc_rom[87] <= 8188;
      adc_rom[88] <= 8185;
      adc_rom[89] <= 8187;
      adc_rom[90] <= 8187;
      adc_rom[91] <= 8183;
      adc_rom[92] <= 8189;
      adc_rom[93] <= 8185;
      adc_rom[94] <= 8188;
      adc_rom[95] <= 8186;
      adc_rom[96] <= 8187;
      adc_rom[97] <= 8189;
      adc_rom[98] <= 8184;
      adc_rom[99] <= 8186;
      adc_rom[100] <= 8185;
      adc_rom[101] <= 8187;
      adc_rom[102] <= 8186;
      adc_rom[103] <= 8184;
      adc_rom[104] <= 8185;
      adc_rom[105] <= 8185;
      adc_rom[106] <= 8187;
      adc_rom[107] <= 8185;
      adc_rom[108] <= 8187;
      adc_rom[109] <= 8185;
      adc_rom[110] <= 8187;
      adc_rom[111] <= 8187;
      adc_rom[112] <= 8188;
      adc_rom[113] <= 8187;
      adc_rom[114] <= 8186;
      adc_rom[115] <= 8187;
      adc_rom[116] <= 8185;
      adc_rom[117] <= 8186;
      adc_rom[118] <= 8184;
      adc_rom[119] <= 8187;
      adc_rom[120] <= 8186;
      adc_rom[121] <= 8186;
      adc_rom[122] <= 8188;
      adc_rom[123] <= 8185;
      adc_rom[124] <= 8186;
      adc_rom[125] <= 8187;
      adc_rom[126] <= 8187;
      adc_rom[127] <= 8187;
      adc_rom[128] <= 8185;
      adc_rom[129] <= 8187;
      adc_rom[130] <= 8185;
      adc_rom[131] <= 8187;
      adc_rom[132] <= 8187;
      adc_rom[133] <= 8185;
      adc_rom[134] <= 8187;
      adc_rom[135] <= 8189;
      adc_rom[136] <= 8188;
      adc_rom[137] <= 8186;
      adc_rom[138] <= 8184;
      adc_rom[139] <= 8186;
      adc_rom[140] <= 8186;
      adc_rom[141] <= 8186;
      adc_rom[142] <= 8189;
      adc_rom[143] <= 8185;
      adc_rom[144] <= 8186;
      adc_rom[145] <= 8186;
      adc_rom[146] <= 8187;
      adc_rom[147] <= 8185;
      adc_rom[148] <= 8187;
      adc_rom[149] <= 8187;
      adc_rom[150] <= 8188;
      adc_rom[151] <= 8188;
      adc_rom[152] <= 8186;
      adc_rom[153] <= 8185;
      adc_rom[154] <= 8187;
      adc_rom[155] <= 8184;
      adc_rom[156] <= 8187;
      adc_rom[157] <= 8187;
      adc_rom[158] <= 8185;
      adc_rom[159] <= 8186;
      adc_rom[160] <= 8187;
      adc_rom[161] <= 8186;
      adc_rom[162] <= 8186;
      adc_rom[163] <= 8186;
      adc_rom[164] <= 8186;
      adc_rom[165] <= 8186;
      adc_rom[166] <= 8186;
      adc_rom[167] <= 8189;
      adc_rom[168] <= 8185;
      adc_rom[169] <= 8185;
      adc_rom[170] <= 8186;
      adc_rom[171] <= 8186;
      adc_rom[172] <= 8186;
      adc_rom[173] <= 8185;
      adc_rom[174] <= 8188;
      adc_rom[175] <= 8185;
      adc_rom[176] <= 8186;
      adc_rom[177] <= 8186;
      adc_rom[178] <= 8187;
      adc_rom[179] <= 8187;
      adc_rom[180] <= 8187;
      adc_rom[181] <= 8187;
      adc_rom[182] <= 8186;
      adc_rom[183] <= 8186;
      adc_rom[184] <= 8187;
      adc_rom[185] <= 8186;
      adc_rom[186] <= 8186;
      adc_rom[187] <= 8187;
      adc_rom[188] <= 8187;
      adc_rom[189] <= 8188;
      adc_rom[190] <= 8185;
      adc_rom[191] <= 8187;
      adc_rom[192] <= 8186;
      adc_rom[193] <= 8187;
      adc_rom[194] <= 8187;
      adc_rom[195] <= 8184;
      adc_rom[196] <= 8187;
      adc_rom[197] <= 8186;
      adc_rom[198] <= 8185;
      adc_rom[199] <= 8187;
      adc_rom[200] <= 8185;
      adc_rom[201] <= 8187;
      adc_rom[202] <= 8185;
      adc_rom[203] <= 8184;
      adc_rom[204] <= 8187;
      adc_rom[205] <= 8185;
      adc_rom[206] <= 8186;
      adc_rom[207] <= 8188;
      adc_rom[208] <= 8185;
      adc_rom[209] <= 8188;
      adc_rom[210] <= 8185;
      adc_rom[211] <= 8187;
      adc_rom[212] <= 8186;
      adc_rom[213] <= 8185;
      adc_rom[214] <= 8184;
      adc_rom[215] <= 8185;
      adc_rom[216] <= 8186;
      adc_rom[217] <= 8186;
      adc_rom[218] <= 8184;
      adc_rom[219] <= 8186;
      adc_rom[220] <= 8185;
      adc_rom[221] <= 8187;
      adc_rom[222] <= 8188;
      adc_rom[223] <= 8185;
      adc_rom[224] <= 8188;
      adc_rom[225] <= 8186;
      adc_rom[226] <= 8186;
      adc_rom[227] <= 8186;
      adc_rom[228] <= 8186;
      adc_rom[229] <= 8189;
      adc_rom[230] <= 8187;
      adc_rom[231] <= 8186;
      adc_rom[232] <= 8187;
      adc_rom[233] <= 8184;
      adc_rom[234] <= 8187;
      adc_rom[235] <= 8187;
      adc_rom[236] <= 8187;
      adc_rom[237] <= 8186;
      adc_rom[238] <= 8185;
      adc_rom[239] <= 8187;
      adc_rom[240] <= 8188;
      adc_rom[241] <= 8185;
      adc_rom[242] <= 8186;
      adc_rom[243] <= 8185;
      adc_rom[244] <= 8186;
      adc_rom[245] <= 8185;
      adc_rom[246] <= 8187;
      adc_rom[247] <= 8187;
      adc_rom[248] <= 8185;
      adc_rom[249] <= 8186;
      adc_rom[250] <= 8185;
      adc_rom[251] <= 8186;
      adc_rom[252] <= 8185;
      adc_rom[253] <= 8185;
      adc_rom[254] <= 8185;
      adc_rom[255] <= 8185;
      adc_rom[256] <= 8187;
      adc_rom[257] <= 8185;
      adc_rom[258] <= 8184;
      adc_rom[259] <= 8186;
      adc_rom[260] <= 8185;
      adc_rom[261] <= 8187;
      adc_rom[262] <= 8186;
      adc_rom[263] <= 8186;
      adc_rom[264] <= 8187;
      adc_rom[265] <= 8186;
      adc_rom[266] <= 8187;
      adc_rom[267] <= 8187;
      adc_rom[268] <= 8186;
      adc_rom[269] <= 8187;
      adc_rom[270] <= 8187;
      adc_rom[271] <= 8187;
      adc_rom[272] <= 8189;
      adc_rom[273] <= 8185;
      adc_rom[274] <= 8188;
      adc_rom[275] <= 8186;
      adc_rom[276] <= 8187;
      adc_rom[277] <= 8187;
      adc_rom[278] <= 8184;
      adc_rom[279] <= 8187;
      adc_rom[280] <= 8187;
      adc_rom[281] <= 8186;
      adc_rom[282] <= 8188;
      adc_rom[283] <= 8187;
      adc_rom[284] <= 8187;
      adc_rom[285] <= 8186;
      adc_rom[286] <= 8186;
      adc_rom[287] <= 8189;
      adc_rom[288] <= 8186;
      adc_rom[289] <= 8186;
      adc_rom[290] <= 8187;
      adc_rom[291] <= 8186;
      adc_rom[292] <= 8185;
      adc_rom[293] <= 8186;
      adc_rom[294] <= 8189;
      adc_rom[295] <= 8185;
      adc_rom[296] <= 8188;
      adc_rom[297] <= 8186;
      adc_rom[298] <= 8186;
      adc_rom[299] <= 8184;
      adc_rom[300] <= 8185;
      adc_rom[301] <= 8185;
      adc_rom[302] <= 8187;
      adc_rom[303] <= 8185;
      adc_rom[304] <= 8185;
      adc_rom[305] <= 8185;
      adc_rom[306] <= 8187;
      adc_rom[307] <= 8184;
      adc_rom[308] <= 8185;
      adc_rom[309] <= 8187;
      adc_rom[310] <= 8186;
      adc_rom[311] <= 8187;
      adc_rom[312] <= 8186;
      adc_rom[313] <= 8184;
      adc_rom[314] <= 8185;
      adc_rom[315] <= 8184;
      adc_rom[316] <= 8185;
      adc_rom[317] <= 8186;
      adc_rom[318] <= 8185;
      adc_rom[319] <= 8187;
      adc_rom[320] <= 8186;
      adc_rom[321] <= 8185;
      adc_rom[322] <= 8186;
      adc_rom[323] <= 8184;
      adc_rom[324] <= 8187;
      adc_rom[325] <= 8186;
      adc_rom[326] <= 8185;
      adc_rom[327] <= 8186;
      adc_rom[328] <= 8182;
      adc_rom[329] <= 8187;
      adc_rom[330] <= 8187;
      adc_rom[331] <= 8186;
      adc_rom[332] <= 8186;
      adc_rom[333] <= 8184;
      adc_rom[334] <= 8183;
      adc_rom[335] <= 8183;
      adc_rom[336] <= 8186;
      adc_rom[337] <= 8185;
      adc_rom[338] <= 8185;
      adc_rom[339] <= 8184;
      adc_rom[340] <= 8186;
      adc_rom[341] <= 8186;
      adc_rom[342] <= 8186;
      adc_rom[343] <= 8185;
      adc_rom[344] <= 8185;
      adc_rom[345] <= 8185;
      adc_rom[346] <= 8183;
      adc_rom[347] <= 8188;
      adc_rom[348] <= 8184;
      adc_rom[349] <= 8187;
      adc_rom[350] <= 8185;
      adc_rom[351] <= 8188;
      adc_rom[352] <= 8186;
      adc_rom[353] <= 8186;
      adc_rom[354] <= 8188;
      adc_rom[355] <= 8184;
      adc_rom[356] <= 8187;
      adc_rom[357] <= 8187;
      adc_rom[358] <= 8185;
      adc_rom[359] <= 8187;
      adc_rom[360] <= 8188;
      adc_rom[361] <= 8187;
      adc_rom[362] <= 8187;
      adc_rom[363] <= 8185;
      adc_rom[364] <= 8188;
      adc_rom[365] <= 8186;
      adc_rom[366] <= 8186;
      adc_rom[367] <= 8186;
      adc_rom[368] <= 8186;
      adc_rom[369] <= 8187;
      adc_rom[370] <= 8187;
      adc_rom[371] <= 8186;
      adc_rom[372] <= 8187;
      adc_rom[373] <= 8185;
      adc_rom[374] <= 8187;
      adc_rom[375] <= 8186;
      adc_rom[376] <= 8186;
      adc_rom[377] <= 8187;
      adc_rom[378] <= 8186;
      adc_rom[379] <= 8190;
      adc_rom[380] <= 8186;
      adc_rom[381] <= 8185;
      adc_rom[382] <= 8187;
      adc_rom[383] <= 8185;
      adc_rom[384] <= 8187;
      adc_rom[385] <= 8186;
      adc_rom[386] <= 8188;
      adc_rom[387] <= 8186;
      adc_rom[388] <= 8186;
      adc_rom[389] <= 8189;
      adc_rom[390] <= 8187;
      adc_rom[391] <= 8188;
      adc_rom[392] <= 8186;
      adc_rom[393] <= 8186;
      adc_rom[394] <= 8188;
      adc_rom[395] <= 8187;
      adc_rom[396] <= 8185;
      adc_rom[397] <= 8187;
      adc_rom[398] <= 8186;
      adc_rom[399] <= 8187;
      adc_rom[400] <= 8187;
      adc_rom[401] <= 8188;
      adc_rom[402] <= 8186;
      adc_rom[403] <= 8185;
      adc_rom[404] <= 8187;
      adc_rom[405] <= 8186;
      adc_rom[406] <= 8186;
      adc_rom[407] <= 8186;
      adc_rom[408] <= 8185;
      adc_rom[409] <= 8186;
      adc_rom[410] <= 8185;
      adc_rom[411] <= 8186;
      adc_rom[412] <= 8187;
      adc_rom[413] <= 8186;
      adc_rom[414] <= 8187;
      adc_rom[415] <= 8185;
      adc_rom[416] <= 8185;
      adc_rom[417] <= 8185;
      adc_rom[418] <= 8184;
      adc_rom[419] <= 8187;
      adc_rom[420] <= 8186;
      adc_rom[421] <= 8186;
      adc_rom[422] <= 8187;
      adc_rom[423] <= 8186;
      adc_rom[424] <= 8187;
      adc_rom[425] <= 8187;
      adc_rom[426] <= 8186;
      adc_rom[427] <= 8186;
      adc_rom[428] <= 8185;
      adc_rom[429] <= 8186;
      adc_rom[430] <= 8185;
      adc_rom[431] <= 8186;
      adc_rom[432] <= 8188;
      adc_rom[433] <= 8184;
      adc_rom[434] <= 8185;
      adc_rom[435] <= 8183;
      adc_rom[436] <= 8189;
      adc_rom[437] <= 8187;
      adc_rom[438] <= 8185;
      adc_rom[439] <= 8186;
      adc_rom[440] <= 8185;
      adc_rom[441] <= 8187;
      adc_rom[442] <= 8188;
      adc_rom[443] <= 8185;
      adc_rom[444] <= 8187;
      adc_rom[445] <= 8184;
      adc_rom[446] <= 8187;
      adc_rom[447] <= 8187;
      adc_rom[448] <= 8183;
      adc_rom[449] <= 8187;
      adc_rom[450] <= 8186;
      adc_rom[451] <= 8186;
      adc_rom[452] <= 8188;
      adc_rom[453] <= 8185;
      adc_rom[454] <= 8188;
      adc_rom[455] <= 8187;
      adc_rom[456] <= 8187;
      adc_rom[457] <= 8186;
      adc_rom[458] <= 8186;
      adc_rom[459] <= 8187;
      adc_rom[460] <= 8185;
      adc_rom[461] <= 8187;
      adc_rom[462] <= 8187;
      adc_rom[463] <= 8185;
      adc_rom[464] <= 8187;
      adc_rom[465] <= 8187;
      adc_rom[466] <= 8188;
      adc_rom[467] <= 8187;
      adc_rom[468] <= 8187;
      adc_rom[469] <= 8187;
      adc_rom[470] <= 8186;
      adc_rom[471] <= 8186;
      adc_rom[472] <= 8186;
      adc_rom[473] <= 8185;
      adc_rom[474] <= 8185;
      adc_rom[475] <= 8185;
      adc_rom[476] <= 8187;
      adc_rom[477] <= 8188;
      adc_rom[478] <= 8187;
      adc_rom[479] <= 8188;
      adc_rom[480] <= 8186;
      adc_rom[481] <= 8185;
      adc_rom[482] <= 8188;
      adc_rom[483] <= 8187;
      adc_rom[484] <= 8186;
      adc_rom[485] <= 8188;
      adc_rom[486] <= 8187;
      adc_rom[487] <= 8187;
      adc_rom[488] <= 8186;
      adc_rom[489] <= 8186;
      adc_rom[490] <= 8185;
      adc_rom[491] <= 8186;
      adc_rom[492] <= 8187;
      adc_rom[493] <= 8186;
      adc_rom[494] <= 8187;
      adc_rom[495] <= 8184;
      adc_rom[496] <= 8186;
      adc_rom[497] <= 8187;
      adc_rom[498] <= 8185;
      adc_rom[499] <= 8187;
      adc_rom[500] <= 8187;
      adc_rom[501] <= 8186;
      adc_rom[502] <= 8186;
      adc_rom[503] <= 8184;
      adc_rom[504] <= 8186;
      adc_rom[505] <= 8186;
      adc_rom[506] <= 8187;
      adc_rom[507] <= 8187;
      adc_rom[508] <= 8185;
      adc_rom[509] <= 8187;
      adc_rom[510] <= 8185;
      adc_rom[511] <= 8185;
      adc_rom[512] <= 8186;
      adc_rom[513] <= 8183;
      adc_rom[514] <= 8187;
      adc_rom[515] <= 8186;
      adc_rom[516] <= 8186;
      adc_rom[517] <= 8189;
      adc_rom[518] <= 8186;
      adc_rom[519] <= 8188;
      adc_rom[520] <= 8186;
      adc_rom[521] <= 8187;
      adc_rom[522] <= 8187;
      adc_rom[523] <= 8185;
      adc_rom[524] <= 8187;
      adc_rom[525] <= 8187;
      adc_rom[526] <= 8188;
      adc_rom[527] <= 8186;
      adc_rom[528] <= 8187;
      adc_rom[529] <= 8186;
      adc_rom[530] <= 8187;
      adc_rom[531] <= 8186;
      adc_rom[532] <= 8186;
      adc_rom[533] <= 8187;
      adc_rom[534] <= 8187;
      adc_rom[535] <= 8186;
      adc_rom[536] <= 8186;
      adc_rom[537] <= 8189;
      adc_rom[538] <= 8185;
      adc_rom[539] <= 8187;
      adc_rom[540] <= 8187;
      adc_rom[541] <= 8187;
      adc_rom[542] <= 8187;
      adc_rom[543] <= 8187;
      adc_rom[544] <= 8188;
      adc_rom[545] <= 8185;
      adc_rom[546] <= 8186;
      adc_rom[547] <= 8187;
      adc_rom[548] <= 8185;
      adc_rom[549] <= 8186;
      adc_rom[550] <= 8185;
      adc_rom[551] <= 8186;
      adc_rom[552] <= 8187;
      adc_rom[553] <= 8187;
      adc_rom[554] <= 8185;
      adc_rom[555] <= 8185;
      adc_rom[556] <= 8185;
      adc_rom[557] <= 8189;
      adc_rom[558] <= 8187;
      adc_rom[559] <= 8187;
      adc_rom[560] <= 8185;
      adc_rom[561] <= 8185;
      adc_rom[562] <= 8187;
      adc_rom[563] <= 8186;
      adc_rom[564] <= 8188;
      adc_rom[565] <= 8186;
      adc_rom[566] <= 8187;
      adc_rom[567] <= 8186;
      adc_rom[568] <= 8185;
      adc_rom[569] <= 8185;
      adc_rom[570] <= 8185;
      adc_rom[571] <= 8187;
      adc_rom[572] <= 8185;
      adc_rom[573] <= 8185;
      adc_rom[574] <= 8187;
      adc_rom[575] <= 8186;
      adc_rom[576] <= 8188;
      adc_rom[577] <= 8188;
      adc_rom[578] <= 8186;
      adc_rom[579] <= 8188;
      adc_rom[580] <= 8185;
      adc_rom[581] <= 8186;
      adc_rom[582] <= 8187;
      adc_rom[583] <= 8184;
      adc_rom[584] <= 8186;
      adc_rom[585] <= 8188;
      adc_rom[586] <= 8186;
      adc_rom[587] <= 8188;
      adc_rom[588] <= 8183;
      adc_rom[589] <= 8187;
      adc_rom[590] <= 8186;
      adc_rom[591] <= 8189;
      adc_rom[592] <= 8187;
      adc_rom[593] <= 8185;
      adc_rom[594] <= 8188;
      adc_rom[595] <= 8186;
      adc_rom[596] <= 8189;
      adc_rom[597] <= 8186;
      adc_rom[598] <= 8187;
      adc_rom[599] <= 8187;
      adc_rom[600] <= 8186;
      adc_rom[601] <= 8187;
      adc_rom[602] <= 8184;
      adc_rom[603] <= 8183;
      adc_rom[604] <= 8188;
      adc_rom[605] <= 8184;
      adc_rom[606] <= 8186;
      adc_rom[607] <= 8185;
      adc_rom[608] <= 8183;
      adc_rom[609] <= 8187;
      adc_rom[610] <= 8186;
      adc_rom[611] <= 8187;
      adc_rom[612] <= 8186;
      adc_rom[613] <= 8185;
      adc_rom[614] <= 8185;
      adc_rom[615] <= 8185;
      adc_rom[616] <= 8185;
      adc_rom[617] <= 8185;
      adc_rom[618] <= 8187;
      adc_rom[619] <= 8188;
      adc_rom[620] <= 8187;
      adc_rom[621] <= 8186;
      adc_rom[622] <= 8187;
      adc_rom[623] <= 8188;
      adc_rom[624] <= 8185;
      adc_rom[625] <= 8185;
      adc_rom[626] <= 8187;
      adc_rom[627] <= 8187;
      adc_rom[628] <= 8185;
      adc_rom[629] <= 8189;
      adc_rom[630] <= 8183;
      adc_rom[631] <= 8186;
      adc_rom[632] <= 8185;
      adc_rom[633] <= 8184;
      adc_rom[634] <= 8186;
      adc_rom[635] <= 8185;
      adc_rom[636] <= 8187;
      adc_rom[637] <= 8186;
      adc_rom[638] <= 8185;
      adc_rom[639] <= 8187;
      adc_rom[640] <= 8186;
      adc_rom[641] <= 8185;
      adc_rom[642] <= 8187;
      adc_rom[643] <= 8186;
      adc_rom[644] <= 8188;
      adc_rom[645] <= 8185;
      adc_rom[646] <= 8185;
      adc_rom[647] <= 8187;
      adc_rom[648] <= 8186;
      adc_rom[649] <= 8185;
      adc_rom[650] <= 8185;
      adc_rom[651] <= 8187;
      adc_rom[652] <= 8186;
      adc_rom[653] <= 8184;
      adc_rom[654] <= 8186;
      adc_rom[655] <= 8184;
      adc_rom[656] <= 8185;
      adc_rom[657] <= 8186;
      adc_rom[658] <= 8185;
      adc_rom[659] <= 8187;
      adc_rom[660] <= 8184;
      adc_rom[661] <= 8185;
      adc_rom[662] <= 8186;
      adc_rom[663] <= 8186;
      adc_rom[664] <= 8186;
      adc_rom[665] <= 8184;
      adc_rom[666] <= 8187;
      adc_rom[667] <= 8185;
      adc_rom[668] <= 8185;
      adc_rom[669] <= 8187;
      adc_rom[670] <= 8185;
      adc_rom[671] <= 8186;
      adc_rom[672] <= 8187;
      adc_rom[673] <= 8185;
      adc_rom[674] <= 8186;
      adc_rom[675] <= 8184;
      adc_rom[676] <= 8186;
      adc_rom[677] <= 8189;
      adc_rom[678] <= 8185;
      adc_rom[679] <= 8184;
      adc_rom[680] <= 8184;
      adc_rom[681] <= 8184;
      adc_rom[682] <= 8184;
      adc_rom[683] <= 8184;
      adc_rom[684] <= 8187;
      adc_rom[685] <= 8182;
      adc_rom[686] <= 8185;
      adc_rom[687] <= 8185;
      adc_rom[688] <= 8184;
      adc_rom[689] <= 8187;
      adc_rom[690] <= 8184;
      adc_rom[691] <= 8185;
      adc_rom[692] <= 8186;
      adc_rom[693] <= 8184;
      adc_rom[694] <= 8186;
      adc_rom[695] <= 8186;
      adc_rom[696] <= 8184;
      adc_rom[697] <= 8187;
      adc_rom[698] <= 8187;
      adc_rom[699] <= 8186;
      adc_rom[700] <= 8185;
      adc_rom[701] <= 8185;
      adc_rom[702] <= 8185;
      adc_rom[703] <= 8184;
      adc_rom[704] <= 8184;
      adc_rom[705] <= 8186;
      adc_rom[706] <= 8184;
      adc_rom[707] <= 8187;
      adc_rom[708] <= 8186;
      adc_rom[709] <= 8189;
      adc_rom[710] <= 8184;
      adc_rom[711] <= 8186;
      adc_rom[712] <= 8184;
      adc_rom[713] <= 8186;
      adc_rom[714] <= 8187;
      adc_rom[715] <= 8186;
      adc_rom[716] <= 8186;
      adc_rom[717] <= 8185;
      adc_rom[718] <= 8186;
      adc_rom[719] <= 8185;
      adc_rom[720] <= 8185;
      adc_rom[721] <= 8185;
      adc_rom[722] <= 8187;
      adc_rom[723] <= 8184;
      adc_rom[724] <= 8186;
      adc_rom[725] <= 8185;
      adc_rom[726] <= 8186;
      adc_rom[727] <= 8187;
      adc_rom[728] <= 8186;
      adc_rom[729] <= 8187;
      adc_rom[730] <= 8184;
      adc_rom[731] <= 8186;
      adc_rom[732] <= 8186;
      adc_rom[733] <= 8186;
      adc_rom[734] <= 8186;
      adc_rom[735] <= 8184;
      adc_rom[736] <= 8187;
      adc_rom[737] <= 8187;
      adc_rom[738] <= 8186;
      adc_rom[739] <= 8183;
      adc_rom[740] <= 8186;
      adc_rom[741] <= 8186;
      adc_rom[742] <= 8186;
      adc_rom[743] <= 8183;
      adc_rom[744] <= 8186;
      adc_rom[745] <= 8186;
      adc_rom[746] <= 8187;
      adc_rom[747] <= 8186;
      adc_rom[748] <= 8183;
      adc_rom[749] <= 8185;
      adc_rom[750] <= 8185;
      adc_rom[751] <= 8185;
      adc_rom[752] <= 8185;
      adc_rom[753] <= 8184;
      adc_rom[754] <= 8187;
      adc_rom[755] <= 8184;
      adc_rom[756] <= 8187;
      adc_rom[757] <= 8186;
      adc_rom[758] <= 8186;
      adc_rom[759] <= 8186;
      adc_rom[760] <= 8186;
      adc_rom[761] <= 8186;
      adc_rom[762] <= 8185;
      adc_rom[763] <= 8186;
      adc_rom[764] <= 8186;
      adc_rom[765] <= 8187;
      adc_rom[766] <= 8184;
      adc_rom[767] <= 8186;
      adc_rom[768] <= 8184;
      adc_rom[769] <= 8188;
      adc_rom[770] <= 8187;
      adc_rom[771] <= 8186;
      adc_rom[772] <= 8186;
      adc_rom[773] <= 8183;
      adc_rom[774] <= 8186;
      adc_rom[775] <= 8184;
      adc_rom[776] <= 8185;
      adc_rom[777] <= 8185;
      adc_rom[778] <= 8184;
      adc_rom[779] <= 8187;
      adc_rom[780] <= 8184;
      adc_rom[781] <= 8187;
      adc_rom[782] <= 8188;
      adc_rom[783] <= 8184;
      adc_rom[784] <= 8186;
      adc_rom[785] <= 8185;
      adc_rom[786] <= 8185;
      adc_rom[787] <= 8186;
      adc_rom[788] <= 8187;
      adc_rom[789] <= 8188;
      adc_rom[790] <= 8185;
      adc_rom[791] <= 8186;
      adc_rom[792] <= 8186;
      adc_rom[793] <= 8186;
      adc_rom[794] <= 8187;
      adc_rom[795] <= 8186;
      adc_rom[796] <= 8186;
      adc_rom[797] <= 8184;
      adc_rom[798] <= 8186;
      adc_rom[799] <= 8188;
      adc_rom[800] <= 8185;
      adc_rom[801] <= 8185;
      adc_rom[802] <= 8186;
      adc_rom[803] <= 8186;
      adc_rom[804] <= 8186;
      adc_rom[805] <= 8186;
      adc_rom[806] <= 8185;
      adc_rom[807] <= 8184;
      adc_rom[808] <= 8184;
      adc_rom[809] <= 8186;
      adc_rom[810] <= 8185;
      adc_rom[811] <= 8188;
      adc_rom[812] <= 8186;
      adc_rom[813] <= 8186;
      adc_rom[814] <= 8189;
      adc_rom[815] <= 8186;
      adc_rom[816] <= 8186;
      adc_rom[817] <= 8187;
      adc_rom[818] <= 8185;
      adc_rom[819] <= 8186;
      adc_rom[820] <= 8186;
      adc_rom[821] <= 8186;
      adc_rom[822] <= 8187;
      adc_rom[823] <= 8186;
      adc_rom[824] <= 8189;
      adc_rom[825] <= 8187;
      adc_rom[826] <= 8186;
      adc_rom[827] <= 8187;
      adc_rom[828] <= 8186;
      adc_rom[829] <= 8187;
      adc_rom[830] <= 8185;
      adc_rom[831] <= 8187;
      adc_rom[832] <= 8185;
      adc_rom[833] <= 8186;
      adc_rom[834] <= 8186;
      adc_rom[835] <= 8185;
      adc_rom[836] <= 8188;
      adc_rom[837] <= 8187;
      adc_rom[838] <= 8184;
      adc_rom[839] <= 8186;
      adc_rom[840] <= 8186;
      adc_rom[841] <= 8189;
      adc_rom[842] <= 8187;
      adc_rom[843] <= 8185;
      adc_rom[844] <= 8185;
      adc_rom[845] <= 8186;
      adc_rom[846] <= 8186;
      adc_rom[847] <= 8184;
      adc_rom[848] <= 8185;
      adc_rom[849] <= 8187;
      adc_rom[850] <= 8185;
      adc_rom[851] <= 8187;
      adc_rom[852] <= 8186;
      adc_rom[853] <= 8186;
      adc_rom[854] <= 8186;
      adc_rom[855] <= 8187;
      adc_rom[856] <= 8186;
      adc_rom[857] <= 8187;
      adc_rom[858] <= 8186;
      adc_rom[859] <= 8188;
      adc_rom[860] <= 8186;
      adc_rom[861] <= 8185;
      adc_rom[862] <= 8188;
      adc_rom[863] <= 8185;
      adc_rom[864] <= 8186;
      adc_rom[865] <= 8185;
      adc_rom[866] <= 8185;
      adc_rom[867] <= 8186;
      adc_rom[868] <= 8184;
      adc_rom[869] <= 8185;
      adc_rom[870] <= 8185;
      adc_rom[871] <= 8187;
      adc_rom[872] <= 8187;
      adc_rom[873] <= 8185;
      adc_rom[874] <= 8185;
      adc_rom[875] <= 8185;
      adc_rom[876] <= 8186;
      adc_rom[877] <= 8185;
      adc_rom[878] <= 8185;
      adc_rom[879] <= 8188;
      adc_rom[880] <= 8185;
      adc_rom[881] <= 8188;
      adc_rom[882] <= 8186;
      adc_rom[883] <= 8186;
      adc_rom[884] <= 8186;
      adc_rom[885] <= 8186;
      adc_rom[886] <= 8187;
      adc_rom[887] <= 8188;
      adc_rom[888] <= 8184;
      adc_rom[889] <= 8185;
      adc_rom[890] <= 8185;
      adc_rom[891] <= 8187;
      adc_rom[892] <= 8186;
      adc_rom[893] <= 8185;
      adc_rom[894] <= 8189;
      adc_rom[895] <= 8186;
      adc_rom[896] <= 8185;
      adc_rom[897] <= 8185;
      adc_rom[898] <= 8185;
      adc_rom[899] <= 8187;
      adc_rom[900] <= 8185;
      adc_rom[901] <= 8186;
      adc_rom[902] <= 8187;
      adc_rom[903] <= 8188;
      adc_rom[904] <= 8187;
      adc_rom[905] <= 8186;
      adc_rom[906] <= 8185;
      adc_rom[907] <= 8185;
      adc_rom[908] <= 8185;
      adc_rom[909] <= 8187;
      adc_rom[910] <= 8185;
      adc_rom[911] <= 8188;
      adc_rom[912] <= 8189;
      adc_rom[913] <= 8185;
      adc_rom[914] <= 8186;
      adc_rom[915] <= 8185;
      adc_rom[916] <= 8184;
      adc_rom[917] <= 8184;
      adc_rom[918] <= 8186;
      adc_rom[919] <= 8185;
      adc_rom[920] <= 8184;
      adc_rom[921] <= 8188;
      adc_rom[922] <= 8185;
      adc_rom[923] <= 8186;
      adc_rom[924] <= 8185;
      adc_rom[925] <= 8183;
      adc_rom[926] <= 8187;
      adc_rom[927] <= 8186;
      adc_rom[928] <= 8185;
      adc_rom[929] <= 8187;
      adc_rom[930] <= 8185;
      adc_rom[931] <= 8185;
      adc_rom[932] <= 8187;
      adc_rom[933] <= 8186;
      adc_rom[934] <= 8185;
      adc_rom[935] <= 8187;
      adc_rom[936] <= 8186;
      adc_rom[937] <= 8187;
      adc_rom[938] <= 8186;
      adc_rom[939] <= 8189;
      adc_rom[940] <= 8186;
      adc_rom[941] <= 8186;
      adc_rom[942] <= 8187;
      adc_rom[943] <= 8186;
      adc_rom[944] <= 8187;
      adc_rom[945] <= 8186;
      adc_rom[946] <= 8189;
      adc_rom[947] <= 8184;
      adc_rom[948] <= 8186;
      adc_rom[949] <= 8190;
      adc_rom[950] <= 8186;
      adc_rom[951] <= 8186;
      adc_rom[952] <= 8187;
      adc_rom[953] <= 8188;
      adc_rom[954] <= 8187;
      adc_rom[955] <= 8187;
      adc_rom[956] <= 8188;
      adc_rom[957] <= 8187;
      adc_rom[958] <= 8187;
      adc_rom[959] <= 8187;
      adc_rom[960] <= 8187;
      adc_rom[961] <= 8184;
      adc_rom[962] <= 8187;
      adc_rom[963] <= 8185;
      adc_rom[964] <= 8189;
      adc_rom[965] <= 8187;
      adc_rom[966] <= 8187;
      adc_rom[967] <= 8186;
      adc_rom[968] <= 8185;
      adc_rom[969] <= 8187;
      adc_rom[970] <= 8186;
      adc_rom[971] <= 8187;
      adc_rom[972] <= 8188;
      adc_rom[973] <= 8184;
      adc_rom[974] <= 8186;
      adc_rom[975] <= 8186;
      adc_rom[976] <= 8184;
      adc_rom[977] <= 8187;
      adc_rom[978] <= 8186;
      adc_rom[979] <= 8187;
      adc_rom[980] <= 8186;
      adc_rom[981] <= 8186;
      adc_rom[982] <= 8184;
      adc_rom[983] <= 8184;
      adc_rom[984] <= 8186;
      adc_rom[985] <= 8186;
      adc_rom[986] <= 8186;
      adc_rom[987] <= 8187;
      adc_rom[988] <= 8185;
      adc_rom[989] <= 8188;
      adc_rom[990] <= 8183;
      adc_rom[991] <= 8184;
      adc_rom[992] <= 8189;
      adc_rom[993] <= 8185;
      adc_rom[994] <= 8186;
      adc_rom[995] <= 8187;
      adc_rom[996] <= 8186;
      adc_rom[997] <= 8187;
      adc_rom[998] <= 8186;
      adc_rom[999] <= 8186;
      adc_rom[1000] <= 8185;
      adc_rom[1001] <= 8186;
      adc_rom[1002] <= 8189;
      adc_rom[1003] <= 8184;
      adc_rom[1004] <= 8185;
      adc_rom[1005] <= 8185;
      adc_rom[1006] <= 8186;
      adc_rom[1007] <= 8185;
      adc_rom[1008] <= 8186;
      adc_rom[1009] <= 8186;
      adc_rom[1010] <= 8185;
      adc_rom[1011] <= 8188;
      adc_rom[1012] <= 8186;
      adc_rom[1013] <= 8184;
      adc_rom[1014] <= 8187;
      adc_rom[1015] <= 8186;
      adc_rom[1016] <= 8187;
      adc_rom[1017] <= 8188;
      adc_rom[1018] <= 8187;
      adc_rom[1019] <= 8187;
      adc_rom[1020] <= 8183;
      adc_rom[1021] <= 8186;
      adc_rom[1022] <= 8186;
      adc_rom[1023] <= 8185;
      adc_rom[1024] <= 8188;
      adc_rom[1025] <= 8187;
      adc_rom[1026] <= 8186;
      adc_rom[1027] <= 8187;
      adc_rom[1028] <= 8185;
      adc_rom[1029] <= 8186;
      adc_rom[1030] <= 8187;
      adc_rom[1031] <= 8187;
      adc_rom[1032] <= 8186;
      adc_rom[1033] <= 8185;
      adc_rom[1034] <= 8187;
      adc_rom[1035] <= 8186;
      adc_rom[1036] <= 8186;
      adc_rom[1037] <= 8184;
      adc_rom[1038] <= 8185;
      adc_rom[1039] <= 8185;
      adc_rom[1040] <= 8187;
      adc_rom[1041] <= 8185;
      adc_rom[1042] <= 8187;
      adc_rom[1043] <= 8185;
      adc_rom[1044] <= 8189;
      adc_rom[1045] <= 8183;
      adc_rom[1046] <= 8187;
      adc_rom[1047] <= 8185;
      adc_rom[1048] <= 8184;
      adc_rom[1049] <= 8186;
      adc_rom[1050] <= 8185;
      adc_rom[1051] <= 8185;
      adc_rom[1052] <= 8189;
      adc_rom[1053] <= 8186;
      adc_rom[1054] <= 8187;
      adc_rom[1055] <= 8185;
      adc_rom[1056] <= 8186;
      adc_rom[1057] <= 8185;
      adc_rom[1058] <= 8187;
      adc_rom[1059] <= 8188;
      adc_rom[1060] <= 8186;
      adc_rom[1061] <= 8186;
      adc_rom[1062] <= 8185;
      adc_rom[1063] <= 8185;
      adc_rom[1064] <= 8188;
      adc_rom[1065] <= 8185;
      adc_rom[1066] <= 8186;
      adc_rom[1067] <= 8186;
      adc_rom[1068] <= 8184;
      adc_rom[1069] <= 8186;
      adc_rom[1070] <= 8186;
      adc_rom[1071] <= 8186;
      adc_rom[1072] <= 8186;
      adc_rom[1073] <= 8184;
      adc_rom[1074] <= 8185;
      adc_rom[1075] <= 8185;
      adc_rom[1076] <= 8186;
      adc_rom[1077] <= 8187;
      adc_rom[1078] <= 8184;
      adc_rom[1079] <= 8186;
      adc_rom[1080] <= 8184;
      adc_rom[1081] <= 8186;
      adc_rom[1082] <= 8187;
      adc_rom[1083] <= 8183;
      adc_rom[1084] <= 8189;
      adc_rom[1085] <= 8185;
      adc_rom[1086] <= 8187;
      adc_rom[1087] <= 8187;
      adc_rom[1088] <= 8184;
      adc_rom[1089] <= 8187;
      adc_rom[1090] <= 8186;
      adc_rom[1091] <= 8186;
      adc_rom[1092] <= 8188;
      adc_rom[1093] <= 8187;
      adc_rom[1094] <= 8189;
      adc_rom[1095] <= 8187;
      adc_rom[1096] <= 8188;
      adc_rom[1097] <= 8186;
      adc_rom[1098] <= 8186;
      adc_rom[1099] <= 8186;
      adc_rom[1100] <= 8187;
      adc_rom[1101] <= 8186;
      adc_rom[1102] <= 8187;
      adc_rom[1103] <= 8184;
      adc_rom[1104] <= 8187;
      adc_rom[1105] <= 8186;
      adc_rom[1106] <= 8187;
      adc_rom[1107] <= 8186;
      adc_rom[1108] <= 8183;
      adc_rom[1109] <= 8187;
      adc_rom[1110] <= 8187;
      adc_rom[1111] <= 8186;
      adc_rom[1112] <= 8186;
      adc_rom[1113] <= 8185;
      adc_rom[1114] <= 8188;
      adc_rom[1115] <= 8185;
      adc_rom[1116] <= 8187;
      adc_rom[1117] <= 8186;
      adc_rom[1118] <= 8187;
      adc_rom[1119] <= 8186;
      adc_rom[1120] <= 8188;
      adc_rom[1121] <= 8186;
      adc_rom[1122] <= 8185;
      adc_rom[1123] <= 8184;
      adc_rom[1124] <= 8187;
      adc_rom[1125] <= 8186;
      adc_rom[1126] <= 8184;
      adc_rom[1127] <= 8187;
      adc_rom[1128] <= 8185;
      adc_rom[1129] <= 8187;
      adc_rom[1130] <= 8187;
      adc_rom[1131] <= 8186;
      adc_rom[1132] <= 8187;
      adc_rom[1133] <= 8184;
      adc_rom[1134] <= 8188;
      adc_rom[1135] <= 8185;
      adc_rom[1136] <= 8186;
      adc_rom[1137] <= 8187;
      adc_rom[1138] <= 8187;
      adc_rom[1139] <= 8187;
      adc_rom[1140] <= 8187;
      adc_rom[1141] <= 8187;
      adc_rom[1142] <= 8189;
      adc_rom[1143] <= 8185;
      adc_rom[1144] <= 8186;
      adc_rom[1145] <= 8184;
      adc_rom[1146] <= 8186;
      adc_rom[1147] <= 8186;
      adc_rom[1148] <= 8187;
      adc_rom[1149] <= 8186;
      adc_rom[1150] <= 8187;
      adc_rom[1151] <= 8186;
      adc_rom[1152] <= 8189;
      adc_rom[1153] <= 8186;
      adc_rom[1154] <= 8186;
      adc_rom[1155] <= 8186;
      adc_rom[1156] <= 8185;
      adc_rom[1157] <= 8186;
      adc_rom[1158] <= 8186;
      adc_rom[1159] <= 8187;
      adc_rom[1160] <= 8183;
      adc_rom[1161] <= 8184;
      adc_rom[1162] <= 8187;
      adc_rom[1163] <= 8186;
      adc_rom[1164] <= 8186;
      adc_rom[1165] <= 8187;
      adc_rom[1166] <= 8187;
      adc_rom[1167] <= 8187;
      adc_rom[1168] <= 8185;
      adc_rom[1169] <= 8186;
      adc_rom[1170] <= 8184;
      adc_rom[1171] <= 8188;
      adc_rom[1172] <= 8187;
      adc_rom[1173] <= 8186;
      adc_rom[1174] <= 8184;
      adc_rom[1175] <= 8186;
      adc_rom[1176] <= 8187;
      adc_rom[1177] <= 8187;
      adc_rom[1178] <= 8185;
      adc_rom[1179] <= 8186;
      adc_rom[1180] <= 8187;
      adc_rom[1181] <= 8187;
      adc_rom[1182] <= 8188;
      adc_rom[1183] <= 8185;
      adc_rom[1184] <= 8186;
      adc_rom[1185] <= 8186;
      adc_rom[1186] <= 8187;
      adc_rom[1187] <= 8186;
      adc_rom[1188] <= 8185;
      adc_rom[1189] <= 8186;
      adc_rom[1190] <= 8185;
      adc_rom[1191] <= 8186;
      adc_rom[1192] <= 8187;
      adc_rom[1193] <= 8184;
      adc_rom[1194] <= 8187;
      adc_rom[1195] <= 8185;
      adc_rom[1196] <= 8186;
      adc_rom[1197] <= 8188;
      adc_rom[1198] <= 8185;
      adc_rom[1199] <= 8187;
      adc_rom[1200] <= 8184;
      adc_rom[1201] <= 8186;
      adc_rom[1202] <= 8188;
      adc_rom[1203] <= 8185;
      adc_rom[1204] <= 8187;
      adc_rom[1205] <= 8185;
      adc_rom[1206] <= 8187;
      adc_rom[1207] <= 8187;
      adc_rom[1208] <= 8185;
      adc_rom[1209] <= 8187;
      adc_rom[1210] <= 8186;
      adc_rom[1211] <= 8187;
      adc_rom[1212] <= 8186;
      adc_rom[1213] <= 8184;
      adc_rom[1214] <= 8186;
      adc_rom[1215] <= 8184;
      adc_rom[1216] <= 8184;
      adc_rom[1217] <= 8186;
      adc_rom[1218] <= 8186;
      adc_rom[1219] <= 8187;
      adc_rom[1220] <= 8184;
      adc_rom[1221] <= 8186;
      adc_rom[1222] <= 8186;
      adc_rom[1223] <= 8185;
      adc_rom[1224] <= 8187;
      adc_rom[1225] <= 8183;
      adc_rom[1226] <= 8187;
      adc_rom[1227] <= 8187;
      adc_rom[1228] <= 8185;
      adc_rom[1229] <= 8187;
      adc_rom[1230] <= 8184;
      adc_rom[1231] <= 8185;
      adc_rom[1232] <= 8185;
      adc_rom[1233] <= 8184;
      adc_rom[1234] <= 8186;
      adc_rom[1235] <= 8185;
      adc_rom[1236] <= 8185;
      adc_rom[1237] <= 8185;
      adc_rom[1238] <= 8183;
      adc_rom[1239] <= 8186;
      adc_rom[1240] <= 8185;
      adc_rom[1241] <= 8185;
      adc_rom[1242] <= 8187;
      adc_rom[1243] <= 8183;
      adc_rom[1244] <= 8185;
      adc_rom[1245] <= 8184;
      adc_rom[1246] <= 8186;
      adc_rom[1247] <= 8187;
      adc_rom[1248] <= 8183;
      adc_rom[1249] <= 8185;
      adc_rom[1250] <= 8187;
      adc_rom[1251] <= 8185;
      adc_rom[1252] <= 8186;
      adc_rom[1253] <= 8186;
      adc_rom[1254] <= 8186;
      adc_rom[1255] <= 8184;
      adc_rom[1256] <= 8186;
      adc_rom[1257] <= 8186;
      adc_rom[1258] <= 8184;
      adc_rom[1259] <= 8184;
      adc_rom[1260] <= 8186;
      adc_rom[1261] <= 8186;
      adc_rom[1262] <= 8187;
      adc_rom[1263] <= 8186;
      adc_rom[1264] <= 8187;
      adc_rom[1265] <= 8186;
      adc_rom[1266] <= 8187;
      adc_rom[1267] <= 8187;
      adc_rom[1268] <= 8184;
      adc_rom[1269] <= 8186;
      adc_rom[1270] <= 8183;
      adc_rom[1271] <= 8187;
      adc_rom[1272] <= 8188;
      adc_rom[1273] <= 8185;
      adc_rom[1274] <= 8189;
      adc_rom[1275] <= 8187;
      adc_rom[1276] <= 8186;
      adc_rom[1277] <= 8188;
      adc_rom[1278] <= 8184;
      adc_rom[1279] <= 8188;
      adc_rom[1280] <= 8186;
      adc_rom[1281] <= 8187;
      adc_rom[1282] <= 8188;
      adc_rom[1283] <= 8184;
      adc_rom[1284] <= 8188;
      adc_rom[1285] <= 8187;
      adc_rom[1286] <= 8186;
      adc_rom[1287] <= 8187;
      adc_rom[1288] <= 8185;
      adc_rom[1289] <= 8188;
      adc_rom[1290] <= 8188;
      adc_rom[1291] <= 8187;
      adc_rom[1292] <= 8186;
      adc_rom[1293] <= 8186;
      adc_rom[1294] <= 8185;
      adc_rom[1295] <= 8184;
      adc_rom[1296] <= 8187;
      adc_rom[1297] <= 8187;
      adc_rom[1298] <= 8184;
      adc_rom[1299] <= 8188;
      adc_rom[1300] <= 8185;
      adc_rom[1301] <= 8184;
      adc_rom[1302] <= 8186;
      adc_rom[1303] <= 8184;
      adc_rom[1304] <= 8187;
      adc_rom[1305] <= 8185;
      adc_rom[1306] <= 8187;
      adc_rom[1307] <= 8187;
      adc_rom[1308] <= 8184;
      adc_rom[1309] <= 8188;
      adc_rom[1310] <= 8184;
      adc_rom[1311] <= 8186;
      adc_rom[1312] <= 8186;
      adc_rom[1313] <= 8184;
      adc_rom[1314] <= 8185;
      adc_rom[1315] <= 8183;
      adc_rom[1316] <= 8185;
      adc_rom[1317] <= 8186;
      adc_rom[1318] <= 8186;
      adc_rom[1319] <= 8186;
      adc_rom[1320] <= 8185;
      adc_rom[1321] <= 8186;
      adc_rom[1322] <= 8187;
      adc_rom[1323] <= 8185;
      adc_rom[1324] <= 8187;
      adc_rom[1325] <= 8186;
      adc_rom[1326] <= 8186;
      adc_rom[1327] <= 8187;
      adc_rom[1328] <= 8186;
      adc_rom[1329] <= 8187;
      adc_rom[1330] <= 8186;
      adc_rom[1331] <= 8186;
      adc_rom[1332] <= 8187;
      adc_rom[1333] <= 8184;
      adc_rom[1334] <= 8186;
      adc_rom[1335] <= 8187;
      adc_rom[1336] <= 8185;
      adc_rom[1337] <= 8188;
      adc_rom[1338] <= 8185;
      adc_rom[1339] <= 8186;
      adc_rom[1340] <= 8186;
      adc_rom[1341] <= 8186;
      adc_rom[1342] <= 8186;
      adc_rom[1343] <= 8186;
      adc_rom[1344] <= 8188;
      adc_rom[1345] <= 8186;
      adc_rom[1346] <= 8186;
      adc_rom[1347] <= 8188;
      adc_rom[1348] <= 8185;
      adc_rom[1349] <= 8185;
      adc_rom[1350] <= 8185;
      adc_rom[1351] <= 8187;
      adc_rom[1352] <= 8187;
      adc_rom[1353] <= 8184;
      adc_rom[1354] <= 8186;
      adc_rom[1355] <= 8183;
      adc_rom[1356] <= 8185;
      adc_rom[1357] <= 8187;
      adc_rom[1358] <= 8185;
      adc_rom[1359] <= 8188;
      adc_rom[1360] <= 8188;
      adc_rom[1361] <= 8186;
      adc_rom[1362] <= 8188;
      adc_rom[1363] <= 8187;
      adc_rom[1364] <= 8186;
      adc_rom[1365] <= 8185;
      adc_rom[1366] <= 8187;
      adc_rom[1367] <= 8184;
      adc_rom[1368] <= 8185;
      adc_rom[1369] <= 8189;
      adc_rom[1370] <= 8187;
      adc_rom[1371] <= 8187;
      adc_rom[1372] <= 8189;
      adc_rom[1373] <= 8185;
      adc_rom[1374] <= 8186;
      adc_rom[1375] <= 8184;
      adc_rom[1376] <= 8187;
      adc_rom[1377] <= 8187;
      adc_rom[1378] <= 8185;
      adc_rom[1379] <= 8188;
      adc_rom[1380] <= 8185;
      adc_rom[1381] <= 8186;
      adc_rom[1382] <= 8184;
      adc_rom[1383] <= 8185;
      adc_rom[1384] <= 8186;
      adc_rom[1385] <= 8185;
      adc_rom[1386] <= 8186;
      adc_rom[1387] <= 8186;
      adc_rom[1388] <= 8186;
      adc_rom[1389] <= 8188;
      adc_rom[1390] <= 8188;
      adc_rom[1391] <= 8188;
      adc_rom[1392] <= 8186;
      adc_rom[1393] <= 8184;
      adc_rom[1394] <= 8186;
      adc_rom[1395] <= 8185;
      adc_rom[1396] <= 8187;
      adc_rom[1397] <= 8187;
      adc_rom[1398] <= 8185;
      adc_rom[1399] <= 8188;
      adc_rom[1400] <= 8185;
      adc_rom[1401] <= 8186;
      adc_rom[1402] <= 8187;
      adc_rom[1403] <= 8185;
      adc_rom[1404] <= 8186;
      adc_rom[1405] <= 8184;
      adc_rom[1406] <= 8189;
      adc_rom[1407] <= 8186;
      adc_rom[1408] <= 8186;
      adc_rom[1409] <= 8186;
      adc_rom[1410] <= 8187;
      adc_rom[1411] <= 8185;
      adc_rom[1412] <= 8188;
      adc_rom[1413] <= 8184;
      adc_rom[1414] <= 8186;
      adc_rom[1415] <= 8185;
      adc_rom[1416] <= 8186;
      adc_rom[1417] <= 8186;
      adc_rom[1418] <= 8185;
      adc_rom[1419] <= 8185;
      adc_rom[1420] <= 8186;
      adc_rom[1421] <= 8186;
      adc_rom[1422] <= 8187;
      adc_rom[1423] <= 8186;
      adc_rom[1424] <= 8188;
      adc_rom[1425] <= 8185;
      adc_rom[1426] <= 8188;
      adc_rom[1427] <= 8189;
      adc_rom[1428] <= 8185;
      adc_rom[1429] <= 8186;
      adc_rom[1430] <= 8184;
      adc_rom[1431] <= 8188;
      adc_rom[1432] <= 8189;
      adc_rom[1433] <= 8185;
      adc_rom[1434] <= 8187;
      adc_rom[1435] <= 8185;
      adc_rom[1436] <= 8185;
      adc_rom[1437] <= 8187;
      adc_rom[1438] <= 8184;
      adc_rom[1439] <= 8189;
      adc_rom[1440] <= 8187;
      adc_rom[1441] <= 8185;
      adc_rom[1442] <= 8185;
      adc_rom[1443] <= 8186;
      adc_rom[1444] <= 8186;
      adc_rom[1445] <= 8185;
      adc_rom[1446] <= 8186;
      adc_rom[1447] <= 8187;
      adc_rom[1448] <= 8188;
      adc_rom[1449] <= 8187;
      adc_rom[1450] <= 8185;
      adc_rom[1451] <= 8187;
      adc_rom[1452] <= 8186;
      adc_rom[1453] <= 8185;
      adc_rom[1454] <= 8187;
      adc_rom[1455] <= 8187;
      adc_rom[1456] <= 8186;
      adc_rom[1457] <= 8186;
      adc_rom[1458] <= 8185;
      adc_rom[1459] <= 8186;
      adc_rom[1460] <= 8185;
      adc_rom[1461] <= 8186;
      adc_rom[1462] <= 8186;
      adc_rom[1463] <= 8184;
      adc_rom[1464] <= 8187;
      adc_rom[1465] <= 8185;
      adc_rom[1466] <= 8186;
      adc_rom[1467] <= 8186;
      adc_rom[1468] <= 8185;
      adc_rom[1469] <= 8187;
      adc_rom[1470] <= 8185;
      adc_rom[1471] <= 8185;
      adc_rom[1472] <= 8186;
      adc_rom[1473] <= 8185;
      adc_rom[1474] <= 8188;
      adc_rom[1475] <= 8185;
      adc_rom[1476] <= 8188;
      adc_rom[1477] <= 8186;
      adc_rom[1478] <= 8185;
      adc_rom[1479] <= 8187;
      adc_rom[1480] <= 8186;
      adc_rom[1481] <= 8186;
      adc_rom[1482] <= 8187;
      adc_rom[1483] <= 8187;
      adc_rom[1484] <= 8188;
      adc_rom[1485] <= 8186;
      adc_rom[1486] <= 8187;
      adc_rom[1487] <= 8187;
      adc_rom[1488] <= 8186;
      adc_rom[1489] <= 8187;
      adc_rom[1490] <= 8186;
      adc_rom[1491] <= 8187;
      adc_rom[1492] <= 8187;
      adc_rom[1493] <= 8188;
      adc_rom[1494] <= 8190;
      adc_rom[1495] <= 8185;
      adc_rom[1496] <= 8186;
      adc_rom[1497] <= 8185;
      adc_rom[1498] <= 8184;
      adc_rom[1499] <= 8187;
      adc_rom[1500] <= 8185;
      adc_rom[1501] <= 8186;
      adc_rom[1502] <= 8187;
      adc_rom[1503] <= 8185;
      adc_rom[1504] <= 8186;
      adc_rom[1505] <= 8186;
      adc_rom[1506] <= 8188;
      adc_rom[1507] <= 8185;
      adc_rom[1508] <= 8185;
      adc_rom[1509] <= 8189;
      adc_rom[1510] <= 8186;
      adc_rom[1511] <= 8185;
      adc_rom[1512] <= 8186;
      adc_rom[1513] <= 8185;
      adc_rom[1514] <= 8188;
      adc_rom[1515] <= 8186;
      adc_rom[1516] <= 8186;
      adc_rom[1517] <= 8187;
      adc_rom[1518] <= 8185;
      adc_rom[1519] <= 8188;
      adc_rom[1520] <= 8186;
      adc_rom[1521] <= 8186;
      adc_rom[1522] <= 8187;
      adc_rom[1523] <= 8185;
      adc_rom[1524] <= 8186;
      adc_rom[1525] <= 8188;
      adc_rom[1526] <= 8185;
      adc_rom[1527] <= 8188;
      adc_rom[1528] <= 8185;
      adc_rom[1529] <= 8185;
      adc_rom[1530] <= 8187;
      adc_rom[1531] <= 8188;
      adc_rom[1532] <= 8188;
      adc_rom[1533] <= 8186;
      adc_rom[1534] <= 8188;
      adc_rom[1535] <= 8184;
      adc_rom[1536] <= 8185;
      adc_rom[1537] <= 8187;
      adc_rom[1538] <= 8187;
      adc_rom[1539] <= 8187;
      adc_rom[1540] <= 8185;
      adc_rom[1541] <= 8185;
      adc_rom[1542] <= 8187;
      adc_rom[1543] <= 8186;
      adc_rom[1544] <= 8188;
      adc_rom[1545] <= 8186;
      adc_rom[1546] <= 8187;
      adc_rom[1547] <= 8185;
      adc_rom[1548] <= 8185;
      adc_rom[1549] <= 8189;
      adc_rom[1550] <= 8185;
      adc_rom[1551] <= 8187;
      adc_rom[1552] <= 8184;
      adc_rom[1553] <= 8185;
      adc_rom[1554] <= 8186;
      adc_rom[1555] <= 8184;
      adc_rom[1556] <= 8186;
      adc_rom[1557] <= 8186;
      adc_rom[1558] <= 8185;
      adc_rom[1559] <= 8187;
      adc_rom[1560] <= 8183;
      adc_rom[1561] <= 8187;
      adc_rom[1562] <= 8188;
      adc_rom[1563] <= 8185;
      adc_rom[1564] <= 8189;
      adc_rom[1565] <= 8185;
      adc_rom[1566] <= 8186;
      adc_rom[1567] <= 8187;
      adc_rom[1568] <= 8186;
      adc_rom[1569] <= 8190;
      adc_rom[1570] <= 8187;
      adc_rom[1571] <= 8188;
      adc_rom[1572] <= 8188;
      adc_rom[1573] <= 8187;
      adc_rom[1574] <= 8189;
      adc_rom[1575] <= 8185;
      adc_rom[1576] <= 8186;
      adc_rom[1577] <= 8184;
      adc_rom[1578] <= 8186;
      adc_rom[1579] <= 8187;
      adc_rom[1580] <= 8185;
      adc_rom[1581] <= 8185;
      adc_rom[1582] <= 8186;
      adc_rom[1583] <= 8185;
      adc_rom[1584] <= 8187;
      adc_rom[1585] <= 8186;
      adc_rom[1586] <= 8183;
      adc_rom[1587] <= 8188;
      adc_rom[1588] <= 8186;
      adc_rom[1589] <= 8186;
      adc_rom[1590] <= 8186;
      adc_rom[1591] <= 8186;
      adc_rom[1592] <= 8186;
      adc_rom[1593] <= 8188;
      adc_rom[1594] <= 8186;
      adc_rom[1595] <= 8184;
      adc_rom[1596] <= 8185;
      adc_rom[1597] <= 8187;
      adc_rom[1598] <= 8185;
      adc_rom[1599] <= 8186;
      adc_rom[1600] <= 8187;
      adc_rom[1601] <= 8185;
      adc_rom[1602] <= 8186;
      adc_rom[1603] <= 8183;
      adc_rom[1604] <= 8187;
      adc_rom[1605] <= 8185;
      adc_rom[1606] <= 8185;
      adc_rom[1607] <= 8188;
      adc_rom[1608] <= 8185;
      adc_rom[1609] <= 8189;
      adc_rom[1610] <= 8185;
      adc_rom[1611] <= 8185;
      adc_rom[1612] <= 8185;
      adc_rom[1613] <= 8185;
      adc_rom[1614] <= 8189;
      adc_rom[1615] <= 8186;
      adc_rom[1616] <= 8186;
      adc_rom[1617] <= 8186;
      adc_rom[1618] <= 8185;
      adc_rom[1619] <= 8187;
      adc_rom[1620] <= 8182;
      adc_rom[1621] <= 8187;
      adc_rom[1622] <= 8186;
      adc_rom[1623] <= 8185;
      adc_rom[1624] <= 8187;
      adc_rom[1625] <= 8186;
      adc_rom[1626] <= 8186;
      adc_rom[1627] <= 8186;
      adc_rom[1628] <= 8187;
      adc_rom[1629] <= 8187;
      adc_rom[1630] <= 8185;
      adc_rom[1631] <= 8187;
      adc_rom[1632] <= 8186;
      adc_rom[1633] <= 8186;
      adc_rom[1634] <= 8188;
      adc_rom[1635] <= 8184;
      adc_rom[1636] <= 8188;
      adc_rom[1637] <= 8185;
      adc_rom[1638] <= 8185;
      adc_rom[1639] <= 8187;
      adc_rom[1640] <= 8185;
      adc_rom[1641] <= 8187;
      adc_rom[1642] <= 8185;
      adc_rom[1643] <= 8186;
      adc_rom[1644] <= 8188;
      adc_rom[1645] <= 8186;
      adc_rom[1646] <= 8188;
      adc_rom[1647] <= 8187;
      adc_rom[1648] <= 8186;
      adc_rom[1649] <= 8186;
      adc_rom[1650] <= 8185;
      adc_rom[1651] <= 8187;
      adc_rom[1652] <= 8186;
      adc_rom[1653] <= 8185;
      adc_rom[1654] <= 8187;
      adc_rom[1655] <= 8186;
      adc_rom[1656] <= 8184;
      adc_rom[1657] <= 8185;
      adc_rom[1658] <= 8186;
      adc_rom[1659] <= 8186;
      adc_rom[1660] <= 8185;
      adc_rom[1661] <= 8187;
      adc_rom[1662] <= 8187;
      adc_rom[1663] <= 8184;
      adc_rom[1664] <= 8185;
      adc_rom[1665] <= 8186;
      adc_rom[1666] <= 8189;
      adc_rom[1667] <= 8189;
      adc_rom[1668] <= 8185;
      adc_rom[1669] <= 8188;
      adc_rom[1670] <= 8184;
      adc_rom[1671] <= 8186;
      adc_rom[1672] <= 8188;
      adc_rom[1673] <= 8186;
      adc_rom[1674] <= 8185;
      adc_rom[1675] <= 8186;
      adc_rom[1676] <= 8184;
      adc_rom[1677] <= 8186;
      adc_rom[1678] <= 8185;
      adc_rom[1679] <= 8187;
      adc_rom[1680] <= 8186;
      adc_rom[1681] <= 8186;
      adc_rom[1682] <= 8187;
      adc_rom[1683] <= 8187;
      adc_rom[1684] <= 8186;
      adc_rom[1685] <= 8184;
      adc_rom[1686] <= 8186;
      adc_rom[1687] <= 8186;
      adc_rom[1688] <= 8186;
      adc_rom[1689] <= 8187;
      adc_rom[1690] <= 8187;
      adc_rom[1691] <= 8186;
      adc_rom[1692] <= 8188;
      adc_rom[1693] <= 8184;
      adc_rom[1694] <= 8187;
      adc_rom[1695] <= 8186;
      adc_rom[1696] <= 8186;
      adc_rom[1697] <= 8185;
      adc_rom[1698] <= 8186;
      adc_rom[1699] <= 8189;
      adc_rom[1700] <= 8186;
      adc_rom[1701] <= 8187;
      adc_rom[1702] <= 8187;
      adc_rom[1703] <= 8185;
      adc_rom[1704] <= 8187;
      adc_rom[1705] <= 8186;
      adc_rom[1706] <= 8186;
      adc_rom[1707] <= 8187;
      adc_rom[1708] <= 8187;
      adc_rom[1709] <= 8187;
      adc_rom[1710] <= 8186;
      adc_rom[1711] <= 8185;
      adc_rom[1712] <= 8189;
      adc_rom[1713] <= 8185;
      adc_rom[1714] <= 8186;
      adc_rom[1715] <= 8186;
      adc_rom[1716] <= 8186;
      adc_rom[1717] <= 8188;
      adc_rom[1718] <= 8186;
      adc_rom[1719] <= 8186;
      adc_rom[1720] <= 8186;
      adc_rom[1721] <= 8187;
      adc_rom[1722] <= 8185;
      adc_rom[1723] <= 8186;
      adc_rom[1724] <= 8186;
      adc_rom[1725] <= 8186;
      adc_rom[1726] <= 8187;
      adc_rom[1727] <= 8186;
      adc_rom[1728] <= 8186;
      adc_rom[1729] <= 8187;
      adc_rom[1730] <= 8189;
      adc_rom[1731] <= 8186;
      adc_rom[1732] <= 8188;
      adc_rom[1733] <= 8186;
      adc_rom[1734] <= 8186;
      adc_rom[1735] <= 8184;
      adc_rom[1736] <= 8187;
      adc_rom[1737] <= 8187;
      adc_rom[1738] <= 8185;
      adc_rom[1739] <= 8188;
      adc_rom[1740] <= 8188;
      adc_rom[1741] <= 8188;
      adc_rom[1742] <= 8186;
      adc_rom[1743] <= 8185;
      adc_rom[1744] <= 8187;
      adc_rom[1745] <= 8186;
      adc_rom[1746] <= 8186;
      adc_rom[1747] <= 8187;
      adc_rom[1748] <= 8184;
      adc_rom[1749] <= 8187;
      adc_rom[1750] <= 8188;
      adc_rom[1751] <= 8186;
      adc_rom[1752] <= 8187;
      adc_rom[1753] <= 8185;
      adc_rom[1754] <= 8185;
      adc_rom[1755] <= 8184;
      adc_rom[1756] <= 8188;
      adc_rom[1757] <= 8187;
      adc_rom[1758] <= 8185;
      adc_rom[1759] <= 8186;
      adc_rom[1760] <= 8186;
      adc_rom[1761] <= 8185;
      adc_rom[1762] <= 8185;
      adc_rom[1763] <= 8186;
      adc_rom[1764] <= 8185;
      adc_rom[1765] <= 8186;
      adc_rom[1766] <= 8185;
      adc_rom[1767] <= 8186;
      adc_rom[1768] <= 8183;
      adc_rom[1769] <= 8184;
      adc_rom[1770] <= 8183;
      adc_rom[1771] <= 8185;
      adc_rom[1772] <= 8186;
      adc_rom[1773] <= 8184;
      adc_rom[1774] <= 8186;
      adc_rom[1775] <= 8185;
      adc_rom[1776] <= 8187;
      adc_rom[1777] <= 8186;
      adc_rom[1778] <= 8183;
      adc_rom[1779] <= 8185;
      adc_rom[1780] <= 8186;
      adc_rom[1781] <= 8186;
      adc_rom[1782] <= 8185;
      adc_rom[1783] <= 8185;
      adc_rom[1784] <= 8188;
      adc_rom[1785] <= 8186;
      adc_rom[1786] <= 8188;
      adc_rom[1787] <= 8187;
      adc_rom[1788] <= 8186;
      adc_rom[1789] <= 8187;
      adc_rom[1790] <= 8185;
      adc_rom[1791] <= 8187;
      adc_rom[1792] <= 8188;
      adc_rom[1793] <= 8183;
      adc_rom[1794] <= 8187;
      adc_rom[1795] <= 8187;
      adc_rom[1796] <= 8186;
      adc_rom[1797] <= 8189;
      adc_rom[1798] <= 8185;
      adc_rom[1799] <= 8187;
      adc_rom[1800] <= 8186;
      adc_rom[1801] <= 8189;
      adc_rom[1802] <= 8186;
      adc_rom[1803] <= 8185;
      adc_rom[1804] <= 8188;
      adc_rom[1805] <= 8185;
      adc_rom[1806] <= 8187;
      adc_rom[1807] <= 8188;
      adc_rom[1808] <= 8186;
      adc_rom[1809] <= 8187;
      adc_rom[1810] <= 8186;
      adc_rom[1811] <= 8186;
      adc_rom[1812] <= 8187;
      adc_rom[1813] <= 8186;
      adc_rom[1814] <= 8189;
      adc_rom[1815] <= 8186;
      adc_rom[1816] <= 8186;
      adc_rom[1817] <= 8187;
      adc_rom[1818] <= 8186;
      adc_rom[1819] <= 8188;
      adc_rom[1820] <= 8185;
      adc_rom[1821] <= 8187;
      adc_rom[1822] <= 8186;
      adc_rom[1823] <= 8185;
      adc_rom[1824] <= 8187;
      adc_rom[1825] <= 8185;
      adc_rom[1826] <= 8187;
      adc_rom[1827] <= 8187;
      adc_rom[1828] <= 8184;
      adc_rom[1829] <= 8186;
      adc_rom[1830] <= 8186;
      adc_rom[1831] <= 8186;
      adc_rom[1832] <= 8185;
      adc_rom[1833] <= 8186;
      adc_rom[1834] <= 8188;
      adc_rom[1835] <= 8184;
      adc_rom[1836] <= 8186;
      adc_rom[1837] <= 8186;
      adc_rom[1838] <= 8185;
      adc_rom[1839] <= 8187;
      adc_rom[1840] <= 8187;
      adc_rom[1841] <= 8186;
      adc_rom[1842] <= 8186;
      adc_rom[1843] <= 8187;
      adc_rom[1844] <= 8187;
      adc_rom[1845] <= 8187;
      adc_rom[1846] <= 8187;
      adc_rom[1847] <= 8188;
      adc_rom[1848] <= 8185;
      adc_rom[1849] <= 8188;
      adc_rom[1850] <= 8185;
      adc_rom[1851] <= 8189;
      adc_rom[1852] <= 8185;
      adc_rom[1853] <= 8187;
      adc_rom[1854] <= 8185;
      adc_rom[1855] <= 8187;
      adc_rom[1856] <= 8186;
      adc_rom[1857] <= 8186;
      adc_rom[1858] <= 8185;
      adc_rom[1859] <= 8186;
      adc_rom[1860] <= 8187;
      adc_rom[1861] <= 8186;
      adc_rom[1862] <= 8187;
      adc_rom[1863] <= 8185;
      adc_rom[1864] <= 8187;
      adc_rom[1865] <= 8185;
      adc_rom[1866] <= 8186;
      adc_rom[1867] <= 8187;
      adc_rom[1868] <= 8184;
      adc_rom[1869] <= 8188;
      adc_rom[1870] <= 8185;
      adc_rom[1871] <= 8185;
      adc_rom[1872] <= 8187;
      adc_rom[1873] <= 8186;
      adc_rom[1874] <= 8187;
      adc_rom[1875] <= 8186;
      adc_rom[1876] <= 8185;
      adc_rom[1877] <= 8187;
      adc_rom[1878] <= 8183;
      adc_rom[1879] <= 8189;
      adc_rom[1880] <= 8185;
      adc_rom[1881] <= 8185;
      adc_rom[1882] <= 8189;
      adc_rom[1883] <= 8184;
      adc_rom[1884] <= 8185;
      adc_rom[1885] <= 8189;
      adc_rom[1886] <= 8187;
      adc_rom[1887] <= 8185;
      adc_rom[1888] <= 8186;
      adc_rom[1889] <= 8189;
      adc_rom[1890] <= 8186;
      adc_rom[1891] <= 8186;
      adc_rom[1892] <= 8186;
      adc_rom[1893] <= 8186;
      adc_rom[1894] <= 8188;
      adc_rom[1895] <= 8186;
      adc_rom[1896] <= 8187;
      adc_rom[1897] <= 8185;
      adc_rom[1898] <= 8184;
      adc_rom[1899] <= 8187;
      adc_rom[1900] <= 8186;
      adc_rom[1901] <= 8186;
      adc_rom[1902] <= 8186;
      adc_rom[1903] <= 8187;
      adc_rom[1904] <= 8185;
      adc_rom[1905] <= 8185;
      adc_rom[1906] <= 8187;
      adc_rom[1907] <= 8189;
      adc_rom[1908] <= 8188;
      adc_rom[1909] <= 8189;
      adc_rom[1910] <= 8186;
      adc_rom[1911] <= 8187;
      adc_rom[1912] <= 8185;
      adc_rom[1913] <= 8187;
      adc_rom[1914] <= 8186;
      adc_rom[1915] <= 8187;
      adc_rom[1916] <= 8187;
      adc_rom[1917] <= 8187;
      adc_rom[1918] <= 8186;
      adc_rom[1919] <= 8187;
      adc_rom[1920] <= 8185;
      adc_rom[1921] <= 8187;
      adc_rom[1922] <= 8185;
      adc_rom[1923] <= 8187;
      adc_rom[1924] <= 8186;
      adc_rom[1925] <= 8186;
      adc_rom[1926] <= 8186;
      adc_rom[1927] <= 8187;
      adc_rom[1928] <= 8186;
      adc_rom[1929] <= 8186;
      adc_rom[1930] <= 8186;
      adc_rom[1931] <= 8187;
      adc_rom[1932] <= 8187;
      adc_rom[1933] <= 8187;
      adc_rom[1934] <= 8187;
      adc_rom[1935] <= 8186;
      adc_rom[1936] <= 8185;
      adc_rom[1937] <= 8189;
      adc_rom[1938] <= 8187;
      adc_rom[1939] <= 8185;
      adc_rom[1940] <= 8186;
      adc_rom[1941] <= 8187;
      adc_rom[1942] <= 8185;
      adc_rom[1943] <= 8186;
      adc_rom[1944] <= 8187;
      adc_rom[1945] <= 8187;
      adc_rom[1946] <= 8189;
      adc_rom[1947] <= 8187;
      adc_rom[1948] <= 8185;
      adc_rom[1949] <= 8186;
      adc_rom[1950] <= 8186;
      adc_rom[1951] <= 8187;
      adc_rom[1952] <= 8187;
      adc_rom[1953] <= 8186;
      adc_rom[1954] <= 8188;
      adc_rom[1955] <= 8184;
      adc_rom[1956] <= 8185;
      adc_rom[1957] <= 8187;
      adc_rom[1958] <= 8187;
      adc_rom[1959] <= 8188;
      adc_rom[1960] <= 8187;
      adc_rom[1961] <= 8186;
      adc_rom[1962] <= 8186;
      adc_rom[1963] <= 8185;
      adc_rom[1964] <= 8187;
      adc_rom[1965] <= 8186;
      adc_rom[1966] <= 8186;
      adc_rom[1967] <= 8187;
      adc_rom[1968] <= 8186;
      adc_rom[1969] <= 8187;
      adc_rom[1970] <= 8187;
      adc_rom[1971] <= 8186;
      adc_rom[1972] <= 8186;
      adc_rom[1973] <= 8185;
      adc_rom[1974] <= 8186;
      adc_rom[1975] <= 8182;
      adc_rom[1976] <= 8185;
      adc_rom[1977] <= 8187;
      adc_rom[1978] <= 8186;
      adc_rom[1979] <= 8187;
      adc_rom[1980] <= 8185;
      adc_rom[1981] <= 8185;
      adc_rom[1982] <= 8187;
      adc_rom[1983] <= 8182;
      adc_rom[1984] <= 8187;
      adc_rom[1985] <= 8185;
      adc_rom[1986] <= 8187;
      adc_rom[1987] <= 8186;
      adc_rom[1988] <= 8188;
      adc_rom[1989] <= 8186;
      adc_rom[1990] <= 8188;
      adc_rom[1991] <= 8188;
      adc_rom[1992] <= 8186;
      adc_rom[1993] <= 8186;
      adc_rom[1994] <= 8186;
      adc_rom[1995] <= 8184;
      adc_rom[1996] <= 8187;
      adc_rom[1997] <= 8186;
      adc_rom[1998] <= 8185;
      adc_rom[1999] <= 8187;
      adc_rom[2000] <= 8183;
      adc_rom[2001] <= 8187;
      adc_rom[2002] <= 8187;
      adc_rom[2003] <= 8185;
      adc_rom[2004] <= 8187;
      adc_rom[2005] <= 8184;
      adc_rom[2006] <= 8186;
      adc_rom[2007] <= 8187;
      adc_rom[2008] <= 8185;
      adc_rom[2009] <= 8187;
      adc_rom[2010] <= 8186;
      adc_rom[2011] <= 8188;
      adc_rom[2012] <= 8189;
      adc_rom[2013] <= 8187;
      adc_rom[2014] <= 8188;
      adc_rom[2015] <= 8185;
      adc_rom[2016] <= 8188;
      adc_rom[2017] <= 8187;
      adc_rom[2018] <= 8184;
      adc_rom[2019] <= 8186;
      adc_rom[2020] <= 8186;
      adc_rom[2021] <= 8186;
      adc_rom[2022] <= 8187;
      adc_rom[2023] <= 8185;
      adc_rom[2024] <= 8188;
      adc_rom[2025] <= 8187;
      adc_rom[2026] <= 8187;
      adc_rom[2027] <= 8185;
      adc_rom[2028] <= 8185;
      adc_rom[2029] <= 8187;
      adc_rom[2030] <= 8186;
      adc_rom[2031] <= 8185;
      adc_rom[2032] <= 8187;
      adc_rom[2033] <= 8186;
      adc_rom[2034] <= 8188;
      adc_rom[2035] <= 8185;
      adc_rom[2036] <= 8189;
      adc_rom[2037] <= 8187;
      adc_rom[2038] <= 8186;
      adc_rom[2039] <= 8187;
      adc_rom[2040] <= 8186;
      adc_rom[2041] <= 8187;
      adc_rom[2042] <= 8186;
      adc_rom[2043] <= 8185;
      adc_rom[2044] <= 8185;
      adc_rom[2045] <= 8186;
      adc_rom[2046] <= 8187;
      adc_rom[2047] <= 8186;
      adc_rom[2048] <= 8185;
      adc_rom[2049] <= 8188;
      adc_rom[2050] <= 8185;
      adc_rom[2051] <= 8186;
      adc_rom[2052] <= 8184;
      adc_rom[2053] <= 8186;
      adc_rom[2054] <= 8187;
      adc_rom[2055] <= 8187;
      adc_rom[2056] <= 8186;
      adc_rom[2057] <= 8186;
      adc_rom[2058] <= 8186;
      adc_rom[2059] <= 8186;
      adc_rom[2060] <= 8184;
      adc_rom[2061] <= 8186;
      adc_rom[2062] <= 8187;
      adc_rom[2063] <= 8185;
      adc_rom[2064] <= 8185;
      adc_rom[2065] <= 8185;
      adc_rom[2066] <= 8185;
      adc_rom[2067] <= 8187;
      adc_rom[2068] <= 8186;
      adc_rom[2069] <= 8186;
      adc_rom[2070] <= 8186;
      adc_rom[2071] <= 8185;
      adc_rom[2072] <= 8187;
      adc_rom[2073] <= 8186;
      adc_rom[2074] <= 8188;
      adc_rom[2075] <= 8185;
      adc_rom[2076] <= 8188;
      adc_rom[2077] <= 8186;
      adc_rom[2078] <= 8184;
      adc_rom[2079] <= 8187;
      adc_rom[2080] <= 8185;
      adc_rom[2081] <= 8190;
      adc_rom[2082] <= 8187;
      adc_rom[2083] <= 8185;
      adc_rom[2084] <= 8189;
      adc_rom[2085] <= 8185;
      adc_rom[2086] <= 8186;
      adc_rom[2087] <= 8186;
      adc_rom[2088] <= 8185;
      adc_rom[2089] <= 8186;
      adc_rom[2090] <= 8188;
      adc_rom[2091] <= 8188;
      adc_rom[2092] <= 8183;
      adc_rom[2093] <= 8186;
      adc_rom[2094] <= 8185;
      adc_rom[2095] <= 8184;
      adc_rom[2096] <= 8186;
      adc_rom[2097] <= 8186;
      adc_rom[2098] <= 8186;
      adc_rom[2099] <= 8186;
      adc_rom[2100] <= 8185;
      adc_rom[2101] <= 8186;
      adc_rom[2102] <= 8186;
      adc_rom[2103] <= 8187;
      adc_rom[2104] <= 8188;
      adc_rom[2105] <= 8186;
      adc_rom[2106] <= 8184;
      adc_rom[2107] <= 8186;
      adc_rom[2108] <= 8183;
      adc_rom[2109] <= 8186;
      adc_rom[2110] <= 8185;
      adc_rom[2111] <= 8186;
      adc_rom[2112] <= 8187;
      adc_rom[2113] <= 8184;
      adc_rom[2114] <= 8186;
      adc_rom[2115] <= 8185;
      adc_rom[2116] <= 8186;
      adc_rom[2117] <= 8187;
      adc_rom[2118] <= 8185;
      adc_rom[2119] <= 8187;
      adc_rom[2120] <= 8187;
      adc_rom[2121] <= 8186;
      adc_rom[2122] <= 8187;
      adc_rom[2123] <= 8188;
      adc_rom[2124] <= 8186;
      adc_rom[2125] <= 8187;
      adc_rom[2126] <= 8186;
      adc_rom[2127] <= 8186;
      adc_rom[2128] <= 8186;
      adc_rom[2129] <= 8190;
      adc_rom[2130] <= 8184;
      adc_rom[2131] <= 8186;
      adc_rom[2132] <= 8186;
      adc_rom[2133] <= 8186;
      adc_rom[2134] <= 8186;
      adc_rom[2135] <= 8187;
      adc_rom[2136] <= 8189;
      adc_rom[2137] <= 8185;
      adc_rom[2138] <= 8185;
      adc_rom[2139] <= 8187;
      adc_rom[2140] <= 8185;
      adc_rom[2141] <= 8186;
      adc_rom[2142] <= 8187;
      adc_rom[2143] <= 8187;
      adc_rom[2144] <= 8185;
      adc_rom[2145] <= 8186;
      adc_rom[2146] <= 8186;
      adc_rom[2147] <= 8187;
      adc_rom[2148] <= 8186;
      adc_rom[2149] <= 8189;
      adc_rom[2150] <= 8187;
      adc_rom[2151] <= 8185;
      adc_rom[2152] <= 8187;
      adc_rom[2153] <= 8187;
      adc_rom[2154] <= 8187;
      adc_rom[2155] <= 8187;
      adc_rom[2156] <= 8188;
      adc_rom[2157] <= 8188;
      adc_rom[2158] <= 8186;
      adc_rom[2159] <= 8187;
      adc_rom[2160] <= 8186;
      adc_rom[2161] <= 8186;
      adc_rom[2162] <= 8187;
      adc_rom[2163] <= 8184;
      adc_rom[2164] <= 8189;
      adc_rom[2165] <= 8187;
      adc_rom[2166] <= 8186;
      adc_rom[2167] <= 8188;
      adc_rom[2168] <= 8185;
      adc_rom[2169] <= 8187;
      adc_rom[2170] <= 8187;
      adc_rom[2171] <= 8186;
      adc_rom[2172] <= 8189;
      adc_rom[2173] <= 8186;
      adc_rom[2174] <= 8186;
      adc_rom[2175] <= 8186;
      adc_rom[2176] <= 8187;
      adc_rom[2177] <= 8187;
      adc_rom[2178] <= 8185;
      adc_rom[2179] <= 8190;
      adc_rom[2180] <= 8187;
      adc_rom[2181] <= 8186;
      adc_rom[2182] <= 8187;
      adc_rom[2183] <= 8186;
      adc_rom[2184] <= 8190;
      adc_rom[2185] <= 8187;
      adc_rom[2186] <= 8186;
      adc_rom[2187] <= 8189;
      adc_rom[2188] <= 8186;
      adc_rom[2189] <= 8188;
      adc_rom[2190] <= 8186;
      adc_rom[2191] <= 8187;
      adc_rom[2192] <= 8186;
      adc_rom[2193] <= 8187;
      adc_rom[2194] <= 8187;
      adc_rom[2195] <= 8186;
      adc_rom[2196] <= 8187;
      adc_rom[2197] <= 8187;
      adc_rom[2198] <= 8187;
      adc_rom[2199] <= 8186;
      adc_rom[2200] <= 8188;
      adc_rom[2201] <= 8188;
      adc_rom[2202] <= 8188;
      adc_rom[2203] <= 8186;
      adc_rom[2204] <= 8188;
      adc_rom[2205] <= 8187;
      adc_rom[2206] <= 8188;
      adc_rom[2207] <= 8187;
      adc_rom[2208] <= 8188;
      adc_rom[2209] <= 8189;
      adc_rom[2210] <= 8186;
      adc_rom[2211] <= 8186;
      adc_rom[2212] <= 8186;
      adc_rom[2213] <= 8185;
      adc_rom[2214] <= 8187;
      adc_rom[2215] <= 8185;
      adc_rom[2216] <= 8187;
      adc_rom[2217] <= 8187;
      adc_rom[2218] <= 8187;
      adc_rom[2219] <= 8188;
      adc_rom[2220] <= 8185;
      adc_rom[2221] <= 8187;
      adc_rom[2222] <= 8189;
      adc_rom[2223] <= 8185;
      adc_rom[2224] <= 8189;
      adc_rom[2225] <= 8188;
      adc_rom[2226] <= 8185;
      adc_rom[2227] <= 8187;
      adc_rom[2228] <= 8185;
      adc_rom[2229] <= 8187;
      adc_rom[2230] <= 8186;
      adc_rom[2231] <= 8186;
      adc_rom[2232] <= 8186;
      adc_rom[2233] <= 8186;
      adc_rom[2234] <= 8185;
      adc_rom[2235] <= 8186;
      adc_rom[2236] <= 8186;
      adc_rom[2237] <= 8186;
      adc_rom[2238] <= 8186;
      adc_rom[2239] <= 8188;
      adc_rom[2240] <= 8185;
      adc_rom[2241] <= 8185;
      adc_rom[2242] <= 8187;
      adc_rom[2243] <= 8188;
      adc_rom[2244] <= 8185;
      adc_rom[2245] <= 8185;
      adc_rom[2246] <= 8185;
      adc_rom[2247] <= 8187;
      adc_rom[2248] <= 8187;
      adc_rom[2249] <= 8186;
      adc_rom[2250] <= 8185;
      adc_rom[2251] <= 8186;
      adc_rom[2252] <= 8186;
      adc_rom[2253] <= 8185;
      adc_rom[2254] <= 8187;
      adc_rom[2255] <= 8187;
      adc_rom[2256] <= 8187;
      adc_rom[2257] <= 8187;
      adc_rom[2258] <= 8186;
      adc_rom[2259] <= 8189;
      adc_rom[2260] <= 8188;
      adc_rom[2261] <= 8188;
      adc_rom[2262] <= 8189;
      adc_rom[2263] <= 8184;
      adc_rom[2264] <= 8188;
      adc_rom[2265] <= 8187;
      adc_rom[2266] <= 8186;
      adc_rom[2267] <= 8187;
      adc_rom[2268] <= 8187;
      adc_rom[2269] <= 8186;
      adc_rom[2270] <= 8186;
      adc_rom[2271] <= 8188;
      adc_rom[2272] <= 8187;
      adc_rom[2273] <= 8187;
      adc_rom[2274] <= 8185;
      adc_rom[2275] <= 8186;
      adc_rom[2276] <= 8187;
      adc_rom[2277] <= 8188;
      adc_rom[2278] <= 8185;
      adc_rom[2279] <= 8187;
      adc_rom[2280] <= 8185;
      adc_rom[2281] <= 8187;
      adc_rom[2282] <= 8188;
      adc_rom[2283] <= 8185;
      adc_rom[2284] <= 8187;
      adc_rom[2285] <= 8186;
      adc_rom[2286] <= 8187;
      adc_rom[2287] <= 8188;
      adc_rom[2288] <= 8185;
      adc_rom[2289] <= 8186;
      adc_rom[2290] <= 8186;
      adc_rom[2291] <= 8186;
      adc_rom[2292] <= 8187;
      adc_rom[2293] <= 8186;
      adc_rom[2294] <= 8187;
      adc_rom[2295] <= 8186;
      adc_rom[2296] <= 8185;
      adc_rom[2297] <= 8188;
      adc_rom[2298] <= 8187;
      adc_rom[2299] <= 8189;
      adc_rom[2300] <= 8187;
      adc_rom[2301] <= 8188;
      adc_rom[2302] <= 8189;
      adc_rom[2303] <= 8185;
      adc_rom[2304] <= 8188;
      adc_rom[2305] <= 8186;
      adc_rom[2306] <= 8188;
      adc_rom[2307] <= 8190;
      adc_rom[2308] <= 8185;
      adc_rom[2309] <= 8187;
      adc_rom[2310] <= 8187;
      adc_rom[2311] <= 8188;
      adc_rom[2312] <= 8187;
      adc_rom[2313] <= 8185;
      adc_rom[2314] <= 8187;
      adc_rom[2315] <= 8186;
      adc_rom[2316] <= 8187;
      adc_rom[2317] <= 8186;
      adc_rom[2318] <= 8185;
      adc_rom[2319] <= 8188;
      adc_rom[2320] <= 8185;
      adc_rom[2321] <= 8189;
      adc_rom[2322] <= 8187;
      adc_rom[2323] <= 8185;
      adc_rom[2324] <= 8186;
      adc_rom[2325] <= 8186;
      adc_rom[2326] <= 8190;
      adc_rom[2327] <= 8186;
      adc_rom[2328] <= 8186;
      adc_rom[2329] <= 8190;
      adc_rom[2330] <= 8184;
      adc_rom[2331] <= 8187;
      adc_rom[2332] <= 8189;
      adc_rom[2333] <= 8185;
      adc_rom[2334] <= 8187;
      adc_rom[2335] <= 8186;
      adc_rom[2336] <= 8186;
      adc_rom[2337] <= 8187;
      adc_rom[2338] <= 8187;
      adc_rom[2339] <= 8187;
      adc_rom[2340] <= 8187;
      adc_rom[2341] <= 8187;
      adc_rom[2342] <= 8186;
      adc_rom[2343] <= 8186;
      adc_rom[2344] <= 8189;
      adc_rom[2345] <= 8189;
      adc_rom[2346] <= 8187;
      adc_rom[2347] <= 8187;
      adc_rom[2348] <= 8185;
      adc_rom[2349] <= 8187;
      adc_rom[2350] <= 8186;
      adc_rom[2351] <= 8187;
      adc_rom[2352] <= 8187;
      adc_rom[2353] <= 8186;
      adc_rom[2354] <= 8186;
      adc_rom[2355] <= 8186;
      adc_rom[2356] <= 8187;
      adc_rom[2357] <= 8186;
      adc_rom[2358] <= 8187;
      adc_rom[2359] <= 8187;
      adc_rom[2360] <= 8185;
      adc_rom[2361] <= 8185;
      adc_rom[2362] <= 8185;
      adc_rom[2363] <= 8185;
      adc_rom[2364] <= 8188;
      adc_rom[2365] <= 8186;
      adc_rom[2366] <= 8189;
      adc_rom[2367] <= 8186;
      adc_rom[2368] <= 8187;
      adc_rom[2369] <= 8188;
      adc_rom[2370] <= 8187;
      adc_rom[2371] <= 8188;
      adc_rom[2372] <= 8188;
      adc_rom[2373] <= 8186;
      adc_rom[2374] <= 8191;
      adc_rom[2375] <= 8185;
      adc_rom[2376] <= 8186;
      adc_rom[2377] <= 8188;
      adc_rom[2378] <= 8186;
      adc_rom[2379] <= 8188;
      adc_rom[2380] <= 8185;
      adc_rom[2381] <= 8186;
      adc_rom[2382] <= 8188;
      adc_rom[2383] <= 8184;
      adc_rom[2384] <= 8186;
      adc_rom[2385] <= 8186;
      adc_rom[2386] <= 8187;
      adc_rom[2387] <= 8187;
      adc_rom[2388] <= 8185;
      adc_rom[2389] <= 8189;
      adc_rom[2390] <= 8187;
      adc_rom[2391] <= 8187;
      adc_rom[2392] <= 8188;
      adc_rom[2393] <= 8187;
      adc_rom[2394] <= 8185;
      adc_rom[2395] <= 8185;
      adc_rom[2396] <= 8187;
      adc_rom[2397] <= 8186;
      adc_rom[2398] <= 8186;
      adc_rom[2399] <= 8188;
      adc_rom[2400] <= 8186;
      adc_rom[2401] <= 8187;
      adc_rom[2402] <= 8187;
      adc_rom[2403] <= 8185;
      adc_rom[2404] <= 8187;
      adc_rom[2405] <= 8187;
      adc_rom[2406] <= 8188;
      adc_rom[2407] <= 8186;
      adc_rom[2408] <= 8185;
      adc_rom[2409] <= 8190;
      adc_rom[2410] <= 8188;
      adc_rom[2411] <= 8186;
      adc_rom[2412] <= 8186;
      adc_rom[2413] <= 8185;
      adc_rom[2414] <= 8189;
      adc_rom[2415] <= 8185;
      adc_rom[2416] <= 8186;
      adc_rom[2417] <= 8187;
      adc_rom[2418] <= 8186;
      adc_rom[2419] <= 8186;
      adc_rom[2420] <= 8187;
      adc_rom[2421] <= 8187;
      adc_rom[2422] <= 8186;
      adc_rom[2423] <= 8187;
      adc_rom[2424] <= 8187;
      adc_rom[2425] <= 8186;
      adc_rom[2426] <= 8187;
      adc_rom[2427] <= 8185;
      adc_rom[2428] <= 8188;
      adc_rom[2429] <= 8187;
      adc_rom[2430] <= 8185;
      adc_rom[2431] <= 8187;
      adc_rom[2432] <= 8187;
      adc_rom[2433] <= 8185;
      adc_rom[2434] <= 8189;
      adc_rom[2435] <= 8188;
      adc_rom[2436] <= 8187;
      adc_rom[2437] <= 8188;
      adc_rom[2438] <= 8187;
      adc_rom[2439] <= 8188;
      adc_rom[2440] <= 8188;
      adc_rom[2441] <= 8184;
      adc_rom[2442] <= 8187;
      adc_rom[2443] <= 8185;
      adc_rom[2444] <= 8190;
      adc_rom[2445] <= 8188;
      adc_rom[2446] <= 8184;
      adc_rom[2447] <= 8186;
      adc_rom[2448] <= 8185;
      adc_rom[2449] <= 8188;
      adc_rom[2450] <= 8186;
      adc_rom[2451] <= 8187;
      adc_rom[2452] <= 8186;
      adc_rom[2453] <= 8185;
      adc_rom[2454] <= 8188;
      adc_rom[2455] <= 8186;
      adc_rom[2456] <= 8187;
      adc_rom[2457] <= 8186;
      adc_rom[2458] <= 8185;
      adc_rom[2459] <= 8188;
      adc_rom[2460] <= 8185;
      adc_rom[2461] <= 8187;
      adc_rom[2462] <= 8185;
      adc_rom[2463] <= 8186;
      adc_rom[2464] <= 8187;
      adc_rom[2465] <= 8183;
      adc_rom[2466] <= 8186;
      adc_rom[2467] <= 8186;
      adc_rom[2468] <= 8187;
      adc_rom[2469] <= 8187;
      adc_rom[2470] <= 8185;
      adc_rom[2471] <= 8186;
      adc_rom[2472] <= 8185;
      adc_rom[2473] <= 8184;
      adc_rom[2474] <= 8189;
      adc_rom[2475] <= 8186;
      adc_rom[2476] <= 8187;
      adc_rom[2477] <= 8187;
      adc_rom[2478] <= 8185;
      adc_rom[2479] <= 8187;
      adc_rom[2480] <= 8187;
      adc_rom[2481] <= 8187;
      adc_rom[2482] <= 8189;
      adc_rom[2483] <= 8186;
      adc_rom[2484] <= 8187;
      adc_rom[2485] <= 8186;
      adc_rom[2486] <= 8187;
      adc_rom[2487] <= 8189;
      adc_rom[2488] <= 8189;
      adc_rom[2489] <= 8187;
      adc_rom[2490] <= 8186;
      adc_rom[2491] <= 8187;
      adc_rom[2492] <= 8188;
      adc_rom[2493] <= 8184;
      adc_rom[2494] <= 8186;
      adc_rom[2495] <= 8185;
      adc_rom[2496] <= 8186;
      adc_rom[2497] <= 8186;
      adc_rom[2498] <= 8186;
      adc_rom[2499] <= 8188;
      adc_rom[2500] <= 8186;
      adc_rom[2501] <= 8187;
      adc_rom[2502] <= 8187;
      adc_rom[2503] <= 8185;
      adc_rom[2504] <= 8186;
      adc_rom[2505] <= 8186;
      adc_rom[2506] <= 8187;
      adc_rom[2507] <= 8186;
      adc_rom[2508] <= 8185;
      adc_rom[2509] <= 8188;
      adc_rom[2510] <= 8187;
      adc_rom[2511] <= 8186;
      adc_rom[2512] <= 8187;
      adc_rom[2513] <= 8185;
      adc_rom[2514] <= 8187;
      adc_rom[2515] <= 8188;
      adc_rom[2516] <= 8186;
      adc_rom[2517] <= 8187;
      adc_rom[2518] <= 8184;
      adc_rom[2519] <= 8187;
      adc_rom[2520] <= 8186;
      adc_rom[2521] <= 8187;
      adc_rom[2522] <= 8188;
      adc_rom[2523] <= 8185;
      adc_rom[2524] <= 8184;
      adc_rom[2525] <= 8187;
      adc_rom[2526] <= 8188;
      adc_rom[2527] <= 8187;
      adc_rom[2528] <= 8186;
      adc_rom[2529] <= 8187;
      adc_rom[2530] <= 8185;
      adc_rom[2531] <= 8186;
      adc_rom[2532] <= 8186;
      adc_rom[2533] <= 8185;
      adc_rom[2534] <= 8188;
      adc_rom[2535] <= 8185;
      adc_rom[2536] <= 8187;
      adc_rom[2537] <= 8188;
      adc_rom[2538] <= 8184;
      adc_rom[2539] <= 8187;
      adc_rom[2540] <= 8186;
      adc_rom[2541] <= 8186;
      adc_rom[2542] <= 8185;
      adc_rom[2543] <= 8186;
      adc_rom[2544] <= 8187;
      adc_rom[2545] <= 8187;
      adc_rom[2546] <= 8187;
      adc_rom[2547] <= 8188;
      adc_rom[2548] <= 8185;
      adc_rom[2549] <= 8186;
      adc_rom[2550] <= 8185;
      adc_rom[2551] <= 8186;
      adc_rom[2552] <= 8187;
      adc_rom[2553] <= 8186;
      adc_rom[2554] <= 8185;
      adc_rom[2555] <= 8186;
      adc_rom[2556] <= 8186;
      adc_rom[2557] <= 8188;
      adc_rom[2558] <= 8187;
      adc_rom[2559] <= 8187;
      adc_rom[2560] <= 8187;
      adc_rom[2561] <= 8189;
      adc_rom[2562] <= 8189;
      adc_rom[2563] <= 8186;
      adc_rom[2564] <= 8187;
      adc_rom[2565] <= 8187;
      adc_rom[2566] <= 8185;
      adc_rom[2567] <= 8187;
      adc_rom[2568] <= 8185;
      adc_rom[2569] <= 8188;
      adc_rom[2570] <= 8187;
      adc_rom[2571] <= 8189;
      adc_rom[2572] <= 8187;
      adc_rom[2573] <= 8187;
      adc_rom[2574] <= 8189;
      adc_rom[2575] <= 8186;
      adc_rom[2576] <= 8187;
      adc_rom[2577] <= 8188;
      adc_rom[2578] <= 8186;
      adc_rom[2579] <= 8186;
      adc_rom[2580] <= 8186;
      adc_rom[2581] <= 8187;
      adc_rom[2582] <= 8188;
      adc_rom[2583] <= 8186;
      adc_rom[2584] <= 8189;
      adc_rom[2585] <= 8186;
      adc_rom[2586] <= 8186;
      adc_rom[2587] <= 8188;
      adc_rom[2588] <= 8185;
      adc_rom[2589] <= 8189;
      adc_rom[2590] <= 8186;
      adc_rom[2591] <= 8189;
      adc_rom[2592] <= 8188;
      adc_rom[2593] <= 8185;
      adc_rom[2594] <= 8187;
      adc_rom[2595] <= 8186;
      adc_rom[2596] <= 8186;
      adc_rom[2597] <= 8187;
      adc_rom[2598] <= 8185;
      adc_rom[2599] <= 8187;
      adc_rom[2600] <= 8189;
      adc_rom[2601] <= 8187;
      adc_rom[2602] <= 8187;
      adc_rom[2603] <= 8185;
      adc_rom[2604] <= 8187;
      adc_rom[2605] <= 8187;
      adc_rom[2606] <= 8187;
      adc_rom[2607] <= 8186;
      adc_rom[2608] <= 8187;
      adc_rom[2609] <= 8190;
      adc_rom[2610] <= 8187;
      adc_rom[2611] <= 8187;
      adc_rom[2612] <= 8187;
      adc_rom[2613] <= 8186;
      adc_rom[2614] <= 8186;
      adc_rom[2615] <= 8186;
      adc_rom[2616] <= 8187;
      adc_rom[2617] <= 8189;
      adc_rom[2618] <= 8186;
      adc_rom[2619] <= 8189;
      adc_rom[2620] <= 8186;
      adc_rom[2621] <= 8186;
      adc_rom[2622] <= 8187;
      adc_rom[2623] <= 8187;
      adc_rom[2624] <= 8190;
      adc_rom[2625] <= 8186;
      adc_rom[2626] <= 8187;
      adc_rom[2627] <= 8188;
      adc_rom[2628] <= 8186;
      adc_rom[2629] <= 8187;
      adc_rom[2630] <= 8186;
      adc_rom[2631] <= 8188;
      adc_rom[2632] <= 8186;
      adc_rom[2633] <= 8187;
      adc_rom[2634] <= 8188;
      adc_rom[2635] <= 8188;
      adc_rom[2636] <= 8189;
      adc_rom[2637] <= 8190;
      adc_rom[2638] <= 8188;
      adc_rom[2639] <= 8188;
      adc_rom[2640] <= 8186;
      adc_rom[2641] <= 8187;
      adc_rom[2642] <= 8188;
      adc_rom[2643] <= 8186;
      adc_rom[2644] <= 8187;
      adc_rom[2645] <= 8187;
      adc_rom[2646] <= 8187;
      adc_rom[2647] <= 8188;
      adc_rom[2648] <= 8186;
      adc_rom[2649] <= 8188;
      adc_rom[2650] <= 8186;
      adc_rom[2651] <= 8187;
      adc_rom[2652] <= 8188;
      adc_rom[2653] <= 8186;
      adc_rom[2654] <= 8186;
      adc_rom[2655] <= 8186;
      adc_rom[2656] <= 8190;
      adc_rom[2657] <= 8187;
      adc_rom[2658] <= 8187;
      adc_rom[2659] <= 8186;
      adc_rom[2660] <= 8187;
      adc_rom[2661] <= 8189;
      adc_rom[2662] <= 8187;
      adc_rom[2663] <= 8185;
      adc_rom[2664] <= 8187;
      adc_rom[2665] <= 8185;
      adc_rom[2666] <= 8187;
      adc_rom[2667] <= 8188;
      adc_rom[2668] <= 8185;
      adc_rom[2669] <= 8187;
      adc_rom[2670] <= 8187;
      adc_rom[2671] <= 8186;
      adc_rom[2672] <= 8189;
      adc_rom[2673] <= 8185;
      adc_rom[2674] <= 8187;
      adc_rom[2675] <= 8187;
      adc_rom[2676] <= 8188;
      adc_rom[2677] <= 8187;
      adc_rom[2678] <= 8187;
      adc_rom[2679] <= 8188;
      adc_rom[2680] <= 8187;
      adc_rom[2681] <= 8184;
      adc_rom[2682] <= 8185;
      adc_rom[2683] <= 8187;
      adc_rom[2684] <= 8189;
      adc_rom[2685] <= 8189;
      adc_rom[2686] <= 8189;
      adc_rom[2687] <= 8187;
      adc_rom[2688] <= 8186;
      adc_rom[2689] <= 8189;
      adc_rom[2690] <= 8186;
      adc_rom[2691] <= 8187;
      adc_rom[2692] <= 8187;
      adc_rom[2693] <= 8185;
      adc_rom[2694] <= 8187;
      adc_rom[2695] <= 8187;
      adc_rom[2696] <= 8187;
      adc_rom[2697] <= 8189;
      adc_rom[2698] <= 8185;
      adc_rom[2699] <= 8187;
      adc_rom[2700] <= 8187;
      adc_rom[2701] <= 8189;
      adc_rom[2702] <= 8189;
      adc_rom[2703] <= 8186;
      adc_rom[2704] <= 8186;
      adc_rom[2705] <= 8187;
      adc_rom[2706] <= 8187;
      adc_rom[2707] <= 8188;
      adc_rom[2708] <= 8184;
      adc_rom[2709] <= 8187;
      adc_rom[2710] <= 8186;
      adc_rom[2711] <= 8186;
      adc_rom[2712] <= 8187;
      adc_rom[2713] <= 8185;
      adc_rom[2714] <= 8187;
      adc_rom[2715] <= 8187;
      adc_rom[2716] <= 8187;
      adc_rom[2717] <= 8187;
      adc_rom[2718] <= 8185;
      adc_rom[2719] <= 8188;
      adc_rom[2720] <= 8189;
      adc_rom[2721] <= 8186;
      adc_rom[2722] <= 8187;
      adc_rom[2723] <= 8187;
      adc_rom[2724] <= 8186;
      adc_rom[2725] <= 8185;
      adc_rom[2726] <= 8186;
      adc_rom[2727] <= 8187;
      adc_rom[2728] <= 8188;
      adc_rom[2729] <= 8188;
      adc_rom[2730] <= 8186;
      adc_rom[2731] <= 8185;
      adc_rom[2732] <= 8188;
      adc_rom[2733] <= 8186;
      adc_rom[2734] <= 8187;
      adc_rom[2735] <= 8185;
      adc_rom[2736] <= 8189;
      adc_rom[2737] <= 8185;
      adc_rom[2738] <= 8186;
      adc_rom[2739] <= 8186;
      adc_rom[2740] <= 8185;
      adc_rom[2741] <= 8186;
      adc_rom[2742] <= 8188;
      adc_rom[2743] <= 8186;
      adc_rom[2744] <= 8187;
      adc_rom[2745] <= 8186;
      adc_rom[2746] <= 8186;
      adc_rom[2747] <= 8187;
      adc_rom[2748] <= 8188;
      adc_rom[2749] <= 8190;
      adc_rom[2750] <= 8186;
      adc_rom[2751] <= 8187;
      adc_rom[2752] <= 8187;
      adc_rom[2753] <= 8186;
      adc_rom[2754] <= 8187;
      adc_rom[2755] <= 8188;
      adc_rom[2756] <= 8187;
      adc_rom[2757] <= 8188;
      adc_rom[2758] <= 8186;
      adc_rom[2759] <= 8189;
      adc_rom[2760] <= 8184;
      adc_rom[2761] <= 8187;
      adc_rom[2762] <= 8187;
      adc_rom[2763] <= 8186;
      adc_rom[2764] <= 8187;
      adc_rom[2765] <= 8184;
      adc_rom[2766] <= 8187;
      adc_rom[2767] <= 8186;
      adc_rom[2768] <= 8187;
      adc_rom[2769] <= 8186;
      adc_rom[2770] <= 8185;
      adc_rom[2771] <= 8188;
      adc_rom[2772] <= 8187;
      adc_rom[2773] <= 8184;
      adc_rom[2774] <= 8187;
      adc_rom[2775] <= 8184;
      adc_rom[2776] <= 8187;
      adc_rom[2777] <= 8187;
      adc_rom[2778] <= 8187;
      adc_rom[2779] <= 8185;
      adc_rom[2780] <= 8186;
      adc_rom[2781] <= 8186;
      adc_rom[2782] <= 8187;
      adc_rom[2783] <= 8185;
      adc_rom[2784] <= 8188;
      adc_rom[2785] <= 8186;
      adc_rom[2786] <= 8188;
      adc_rom[2787] <= 8189;
      adc_rom[2788] <= 8186;
      adc_rom[2789] <= 8187;
      adc_rom[2790] <= 8186;
      adc_rom[2791] <= 8187;
      adc_rom[2792] <= 8187;
      adc_rom[2793] <= 8186;
      adc_rom[2794] <= 8187;
      adc_rom[2795] <= 8186;
      adc_rom[2796] <= 8186;
      adc_rom[2797] <= 8186;
      adc_rom[2798] <= 8185;
      adc_rom[2799] <= 8188;
      adc_rom[2800] <= 8186;
      adc_rom[2801] <= 8186;
      adc_rom[2802] <= 8186;
      adc_rom[2803] <= 8184;
      adc_rom[2804] <= 8187;
      adc_rom[2805] <= 8188;
      adc_rom[2806] <= 8186;
      adc_rom[2807] <= 8188;
      adc_rom[2808] <= 8186;
      adc_rom[2809] <= 8186;
      adc_rom[2810] <= 8185;
      adc_rom[2811] <= 8185;
      adc_rom[2812] <= 8186;
      adc_rom[2813] <= 8184;
      adc_rom[2814] <= 8186;
      adc_rom[2815] <= 8185;
      adc_rom[2816] <= 8185;
      adc_rom[2817] <= 8189;
      adc_rom[2818] <= 8185;
      adc_rom[2819] <= 8187;
      adc_rom[2820] <= 8184;
      adc_rom[2821] <= 8187;
      adc_rom[2822] <= 8186;
      adc_rom[2823] <= 8187;
      adc_rom[2824] <= 8187;
      adc_rom[2825] <= 8185;
      adc_rom[2826] <= 8188;
      adc_rom[2827] <= 8188;
      adc_rom[2828] <= 8186;
      adc_rom[2829] <= 8187;
      adc_rom[2830] <= 8183;
      adc_rom[2831] <= 8187;
      adc_rom[2832] <= 8188;
      adc_rom[2833] <= 8185;
      adc_rom[2834] <= 8186;
      adc_rom[2835] <= 8185;
      adc_rom[2836] <= 8186;
      adc_rom[2837] <= 8187;
      adc_rom[2838] <= 8187;
      adc_rom[2839] <= 8188;
      adc_rom[2840] <= 8185;
      adc_rom[2841] <= 8186;
      adc_rom[2842] <= 8186;
      adc_rom[2843] <= 8186;
      adc_rom[2844] <= 8189;
      adc_rom[2845] <= 8187;
      adc_rom[2846] <= 8186;
      adc_rom[2847] <= 8186;
      adc_rom[2848] <= 8186;
      adc_rom[2849] <= 8186;
      adc_rom[2850] <= 8186;
      adc_rom[2851] <= 8186;
      adc_rom[2852] <= 8189;
      adc_rom[2853] <= 8187;
      adc_rom[2854] <= 8188;
      adc_rom[2855] <= 8185;
      adc_rom[2856] <= 8188;
      adc_rom[2857] <= 8188;
      adc_rom[2858] <= 8186;
      adc_rom[2859] <= 8187;
      adc_rom[2860] <= 8187;
      adc_rom[2861] <= 8188;
      adc_rom[2862] <= 8187;
      adc_rom[2863] <= 8187;
      adc_rom[2864] <= 8189;
      adc_rom[2865] <= 8184;
      adc_rom[2866] <= 8186;
      adc_rom[2867] <= 8186;
      adc_rom[2868] <= 8186;
      adc_rom[2869] <= 8189;
      adc_rom[2870] <= 8184;
      adc_rom[2871] <= 8187;
      adc_rom[2872] <= 8186;
      adc_rom[2873] <= 8187;
      adc_rom[2874] <= 8188;
      adc_rom[2875] <= 8187;
      adc_rom[2876] <= 8187;
      adc_rom[2877] <= 8186;
      adc_rom[2878] <= 8186;
      adc_rom[2879] <= 8187;
      adc_rom[2880] <= 8186;
      adc_rom[2881] <= 8187;
      adc_rom[2882] <= 8187;
      adc_rom[2883] <= 8188;
      adc_rom[2884] <= 8189;
      adc_rom[2885] <= 8185;
      adc_rom[2886] <= 8189;
      adc_rom[2887] <= 8188;
      adc_rom[2888] <= 8188;
      adc_rom[2889] <= 8187;
      adc_rom[2890] <= 8186;
      adc_rom[2891] <= 8188;
      adc_rom[2892] <= 8186;
      adc_rom[2893] <= 8186;
      adc_rom[2894] <= 8188;
      adc_rom[2895] <= 8186;
      adc_rom[2896] <= 8187;
      adc_rom[2897] <= 8186;
      adc_rom[2898] <= 8186;
      adc_rom[2899] <= 8187;
      adc_rom[2900] <= 8187;
      adc_rom[2901] <= 8186;
      adc_rom[2902] <= 8186;
      adc_rom[2903] <= 8185;
      adc_rom[2904] <= 8189;
      adc_rom[2905] <= 8186;
      adc_rom[2906] <= 8186;
      adc_rom[2907] <= 8188;
      adc_rom[2908] <= 8185;
      adc_rom[2909] <= 8187;
      adc_rom[2910] <= 8185;
      adc_rom[2911] <= 8186;
      adc_rom[2912] <= 8187;
      adc_rom[2913] <= 8185;
      adc_rom[2914] <= 8188;
      adc_rom[2915] <= 8187;
      adc_rom[2916] <= 8186;
      adc_rom[2917] <= 8187;
      adc_rom[2918] <= 8185;
      adc_rom[2919] <= 8188;
      adc_rom[2920] <= 8187;
      adc_rom[2921] <= 8186;
      adc_rom[2922] <= 8187;
      adc_rom[2923] <= 8186;
      adc_rom[2924] <= 8187;
      adc_rom[2925] <= 8185;
      adc_rom[2926] <= 8185;
      adc_rom[2927] <= 8185;
      adc_rom[2928] <= 8186;
      adc_rom[2929] <= 8188;
      adc_rom[2930] <= 8186;
      adc_rom[2931] <= 8189;
      adc_rom[2932] <= 8189;
      adc_rom[2933] <= 8185;
      adc_rom[2934] <= 8186;
      adc_rom[2935] <= 8186;
      adc_rom[2936] <= 8187;
      adc_rom[2937] <= 8186;
      adc_rom[2938] <= 8185;
      adc_rom[2939] <= 8187;
      adc_rom[2940] <= 8185;
      adc_rom[2941] <= 8186;
      adc_rom[2942] <= 8186;
      adc_rom[2943] <= 8186;
      adc_rom[2944] <= 8186;
      adc_rom[2945] <= 8186;
      adc_rom[2946] <= 8186;
      adc_rom[2947] <= 8187;
      adc_rom[2948] <= 8186;
      adc_rom[2949] <= 8185;
      adc_rom[2950] <= 8186;
      adc_rom[2951] <= 8187;
      adc_rom[2952] <= 8188;
      adc_rom[2953] <= 8185;
      adc_rom[2954] <= 8187;
      adc_rom[2955] <= 8187;
      adc_rom[2956] <= 8184;
      adc_rom[2957] <= 8187;
      adc_rom[2958] <= 8184;
      adc_rom[2959] <= 8189;
      adc_rom[2960] <= 8187;
      adc_rom[2961] <= 8188;
      adc_rom[2962] <= 8189;
      adc_rom[2963] <= 8187;
      adc_rom[2964] <= 8187;
      adc_rom[2965] <= 8184;
      adc_rom[2966] <= 8187;
      adc_rom[2967] <= 8187;
      adc_rom[2968] <= 8185;
      adc_rom[2969] <= 8186;
      adc_rom[2970] <= 8185;
      adc_rom[2971] <= 8186;
      adc_rom[2972] <= 8187;
      adc_rom[2973] <= 8186;
      adc_rom[2974] <= 8186;
      adc_rom[2975] <= 8185;
      adc_rom[2976] <= 8186;
      adc_rom[2977] <= 8187;
      adc_rom[2978] <= 8187;
      adc_rom[2979] <= 8189;
      adc_rom[2980] <= 8185;
      adc_rom[2981] <= 8186;
      adc_rom[2982] <= 8186;
      adc_rom[2983] <= 8186;
      adc_rom[2984] <= 8186;
      adc_rom[2985] <= 8184;
      adc_rom[2986] <= 8186;
      adc_rom[2987] <= 8185;
      adc_rom[2988] <= 8186;
      adc_rom[2989] <= 8187;
      adc_rom[2990] <= 8185;
      adc_rom[2991] <= 8186;
      adc_rom[2992] <= 8186;
      adc_rom[2993] <= 8186;
      adc_rom[2994] <= 8188;
      adc_rom[2995] <= 8186;
      adc_rom[2996] <= 8185;
      adc_rom[2997] <= 8187;
      adc_rom[2998] <= 8186;
      adc_rom[2999] <= 8190;
      adc_rom[3000] <= 8186;
      adc_rom[3001] <= 8187;
      adc_rom[3002] <= 8189;
      adc_rom[3003] <= 8185;
      adc_rom[3004] <= 8188;
      adc_rom[3005] <= 8185;
      adc_rom[3006] <= 8187;
      adc_rom[3007] <= 8186;
      adc_rom[3008] <= 8185;
      adc_rom[3009] <= 8189;
      adc_rom[3010] <= 8186;
      adc_rom[3011] <= 8186;
      adc_rom[3012] <= 8184;
      adc_rom[3013] <= 8187;
      adc_rom[3014] <= 8186;
      adc_rom[3015] <= 8186;
      adc_rom[3016] <= 8185;
      adc_rom[3017] <= 8189;
      adc_rom[3018] <= 8185;
      adc_rom[3019] <= 8187;
      adc_rom[3020] <= 8185;
      adc_rom[3021] <= 8186;
      adc_rom[3022] <= 8187;
      adc_rom[3023] <= 8186;
      adc_rom[3024] <= 8186;
      adc_rom[3025] <= 8186;
      adc_rom[3026] <= 8187;
      adc_rom[3027] <= 8187;
      adc_rom[3028] <= 8186;
      adc_rom[3029] <= 8185;
      adc_rom[3030] <= 8186;
      adc_rom[3031] <= 8187;
      adc_rom[3032] <= 8187;
      adc_rom[3033] <= 8187;
      adc_rom[3034] <= 8186;
      adc_rom[3035] <= 8187;
      adc_rom[3036] <= 8187;
      adc_rom[3037] <= 8188;
      adc_rom[3038] <= 8186;
      adc_rom[3039] <= 8188;
      adc_rom[3040] <= 8187;
      adc_rom[3041] <= 8187;
      adc_rom[3042] <= 8187;
      adc_rom[3043] <= 8182;
      adc_rom[3044] <= 8187;
      adc_rom[3045] <= 8185;
      adc_rom[3046] <= 8186;
      adc_rom[3047] <= 8188;
      adc_rom[3048] <= 8187;
      adc_rom[3049] <= 8188;
      adc_rom[3050] <= 8187;
      adc_rom[3051] <= 8188;
      adc_rom[3052] <= 8186;
      adc_rom[3053] <= 8186;
      adc_rom[3054] <= 8187;
      adc_rom[3055] <= 8187;
      adc_rom[3056] <= 8186;
      adc_rom[3057] <= 8188;
      adc_rom[3058] <= 8186;
      adc_rom[3059] <= 8189;
      adc_rom[3060] <= 8185;
      adc_rom[3061] <= 8189;
      adc_rom[3062] <= 8186;
      adc_rom[3063] <= 8186;
      adc_rom[3064] <= 8185;
      adc_rom[3065] <= 8185;
      adc_rom[3066] <= 8184;
      adc_rom[3067] <= 8186;
      adc_rom[3068] <= 8186;
      adc_rom[3069] <= 8188;
      adc_rom[3070] <= 8186;
      adc_rom[3071] <= 8185;
      adc_rom[3072] <= 8187;
      adc_rom[3073] <= 8184;
      adc_rom[3074] <= 8190;
      adc_rom[3075] <= 8188;
      adc_rom[3076] <= 8186;
      adc_rom[3077] <= 8188;
      adc_rom[3078] <= 8186;
      adc_rom[3079] <= 8190;
      adc_rom[3080] <= 8186;
      adc_rom[3081] <= 8185;
      adc_rom[3082] <= 8187;
      adc_rom[3083] <= 8183;
      adc_rom[3084] <= 8188;
      adc_rom[3085] <= 8186;
      adc_rom[3086] <= 8185;
      adc_rom[3087] <= 8187;
      adc_rom[3088] <= 8185;
      adc_rom[3089] <= 8187;
      adc_rom[3090] <= 8185;
      adc_rom[3091] <= 8185;
      adc_rom[3092] <= 8189;
      adc_rom[3093] <= 8186;
      adc_rom[3094] <= 8188;
      adc_rom[3095] <= 8185;
      adc_rom[3096] <= 8187;
      adc_rom[3097] <= 8187;
      adc_rom[3098] <= 8184;
      adc_rom[3099] <= 8187;
      adc_rom[3100] <= 8185;
      adc_rom[3101] <= 8186;
      adc_rom[3102] <= 8186;
      adc_rom[3103] <= 8186;
      adc_rom[3104] <= 8186;
      adc_rom[3105] <= 8187;
      adc_rom[3106] <= 8185;
      adc_rom[3107] <= 8188;
      adc_rom[3108] <= 8186;
      adc_rom[3109] <= 8186;
      adc_rom[3110] <= 8185;
      adc_rom[3111] <= 8187;
      adc_rom[3112] <= 8186;
      adc_rom[3113] <= 8186;
      adc_rom[3114] <= 8187;
      adc_rom[3115] <= 8185;
      adc_rom[3116] <= 8186;
      adc_rom[3117] <= 8187;
      adc_rom[3118] <= 8187;
      adc_rom[3119] <= 8186;
      adc_rom[3120] <= 8186;
      adc_rom[3121] <= 8187;
      adc_rom[3122] <= 8186;
      adc_rom[3123] <= 8185;
      adc_rom[3124] <= 8187;
      adc_rom[3125] <= 8186;
      adc_rom[3126] <= 8186;
      adc_rom[3127] <= 8186;
      adc_rom[3128] <= 8185;
      adc_rom[3129] <= 8185;
      adc_rom[3130] <= 8186;
      adc_rom[3131] <= 8187;
      adc_rom[3132] <= 8187;
      adc_rom[3133] <= 8184;
      adc_rom[3134] <= 8185;
      adc_rom[3135] <= 8187;
      adc_rom[3136] <= 8187;
      adc_rom[3137] <= 8189;
      adc_rom[3138] <= 8187;
      adc_rom[3139] <= 8187;
      adc_rom[3140] <= 8185;
      adc_rom[3141] <= 8186;
      adc_rom[3142] <= 8186;
      adc_rom[3143] <= 8188;
      adc_rom[3144] <= 8186;
      adc_rom[3145] <= 8186;
      adc_rom[3146] <= 8189;
      adc_rom[3147] <= 8189;
      adc_rom[3148] <= 8185;
      adc_rom[3149] <= 8188;
      adc_rom[3150] <= 8188;
      adc_rom[3151] <= 8187;
      adc_rom[3152] <= 8186;
      adc_rom[3153] <= 8185;
      adc_rom[3154] <= 8186;
      adc_rom[3155] <= 8186;
      adc_rom[3156] <= 8185;
      adc_rom[3157] <= 8188;
      adc_rom[3158] <= 8184;
      adc_rom[3159] <= 8186;
      adc_rom[3160] <= 8185;
      adc_rom[3161] <= 8187;
      adc_rom[3162] <= 8187;
      adc_rom[3163] <= 8184;
      adc_rom[3164] <= 8187;
      adc_rom[3165] <= 8187;
      adc_rom[3166] <= 8190;
      adc_rom[3167] <= 8189;
      adc_rom[3168] <= 8185;
      adc_rom[3169] <= 8188;
      adc_rom[3170] <= 8185;
      adc_rom[3171] <= 8187;
      adc_rom[3172] <= 8185;
      adc_rom[3173] <= 8184;
      adc_rom[3174] <= 8186;
      adc_rom[3175] <= 8187;
      adc_rom[3176] <= 8186;
      adc_rom[3177] <= 8185;
      adc_rom[3178] <= 8186;
      adc_rom[3179] <= 8188;
      adc_rom[3180] <= 8186;
      adc_rom[3181] <= 8186;
      adc_rom[3182] <= 8185;
      adc_rom[3183] <= 8186;
      adc_rom[3184] <= 8187;
      adc_rom[3185] <= 8184;
      adc_rom[3186] <= 8185;
      adc_rom[3187] <= 8188;
      adc_rom[3188] <= 8187;
      adc_rom[3189] <= 8186;
      adc_rom[3190] <= 8185;
      adc_rom[3191] <= 8187;
      adc_rom[3192] <= 8186;
      adc_rom[3193] <= 8184;
      adc_rom[3194] <= 8187;
      adc_rom[3195] <= 8185;
      adc_rom[3196] <= 8185;
      adc_rom[3197] <= 8186;
      adc_rom[3198] <= 8184;
      adc_rom[3199] <= 8186;
      adc_rom[3200] <= 8184;
      adc_rom[3201] <= 8186;
      adc_rom[3202] <= 8187;
      adc_rom[3203] <= 8185;
      adc_rom[3204] <= 8187;
      adc_rom[3205] <= 8187;
      adc_rom[3206] <= 8186;
      adc_rom[3207] <= 8189;
      adc_rom[3208] <= 8185;
      adc_rom[3209] <= 8188;
      adc_rom[3210] <= 8184;
      adc_rom[3211] <= 8186;
      adc_rom[3212] <= 8186;
      adc_rom[3213] <= 8187;
      adc_rom[3214] <= 8188;
      adc_rom[3215] <= 8187;
      adc_rom[3216] <= 8186;
      adc_rom[3217] <= 8187;
      adc_rom[3218] <= 8186;
      adc_rom[3219] <= 8186;
      adc_rom[3220] <= 8188;
      adc_rom[3221] <= 8185;
      adc_rom[3222] <= 8186;
      adc_rom[3223] <= 8186;
      adc_rom[3224] <= 8188;
      adc_rom[3225] <= 8187;
      adc_rom[3226] <= 8186;
      adc_rom[3227] <= 8188;
      adc_rom[3228] <= 8184;
      adc_rom[3229] <= 8184;
      adc_rom[3230] <= 8187;
      adc_rom[3231] <= 8187;
      adc_rom[3232] <= 8188;
      adc_rom[3233] <= 8183;
      adc_rom[3234] <= 8186;
      adc_rom[3235] <= 8183;
      adc_rom[3236] <= 8186;
      adc_rom[3237] <= 8185;
      adc_rom[3238] <= 8185;
      adc_rom[3239] <= 8186;
      adc_rom[3240] <= 8185;
      adc_rom[3241] <= 8188;
      adc_rom[3242] <= 8187;
      adc_rom[3243] <= 8185;
      adc_rom[3244] <= 8187;
      adc_rom[3245] <= 8186;
      adc_rom[3246] <= 8187;
      adc_rom[3247] <= 8187;
      adc_rom[3248] <= 8188;
      adc_rom[3249] <= 8188;
      adc_rom[3250] <= 8186;
      adc_rom[3251] <= 8187;
      adc_rom[3252] <= 8185;
      adc_rom[3253] <= 8185;
      adc_rom[3254] <= 8186;
      adc_rom[3255] <= 8185;
      adc_rom[3256] <= 8186;
      adc_rom[3257] <= 8186;
      adc_rom[3258] <= 8185;
      adc_rom[3259] <= 8187;
      adc_rom[3260] <= 8184;
      adc_rom[3261] <= 8186;
      adc_rom[3262] <= 8186;
      adc_rom[3263] <= 8184;
      adc_rom[3264] <= 8187;
      adc_rom[3265] <= 8185;
      adc_rom[3266] <= 8188;
      adc_rom[3267] <= 8187;
      adc_rom[3268] <= 8185;
      adc_rom[3269] <= 8186;
      adc_rom[3270] <= 8186;
      adc_rom[3271] <= 8186;
      adc_rom[3272] <= 8187;
      adc_rom[3273] <= 8183;
      adc_rom[3274] <= 8185;
      adc_rom[3275] <= 8185;
      adc_rom[3276] <= 8187;
      adc_rom[3277] <= 8185;
      adc_rom[3278] <= 8184;
      adc_rom[3279] <= 8187;
      adc_rom[3280] <= 8187;
      adc_rom[3281] <= 8188;
      adc_rom[3282] <= 8187;
      adc_rom[3283] <= 8184;
      adc_rom[3284] <= 8187;
      adc_rom[3285] <= 8186;
      adc_rom[3286] <= 8187;
      adc_rom[3287] <= 8187;
      adc_rom[3288] <= 8186;
      adc_rom[3289] <= 8187;
      adc_rom[3290] <= 8183;
      adc_rom[3291] <= 8187;
      adc_rom[3292] <= 8186;
      adc_rom[3293] <= 8186;
      adc_rom[3294] <= 8187;
      adc_rom[3295] <= 8186;
      adc_rom[3296] <= 8187;
      adc_rom[3297] <= 8185;
      adc_rom[3298] <= 8185;
      adc_rom[3299] <= 8186;
      adc_rom[3300] <= 8186;
      adc_rom[3301] <= 8186;
      adc_rom[3302] <= 8186;
      adc_rom[3303] <= 8186;
      adc_rom[3304] <= 8186;
      adc_rom[3305] <= 8185;
      adc_rom[3306] <= 8185;
      adc_rom[3307] <= 8187;
      adc_rom[3308] <= 8186;
      adc_rom[3309] <= 8185;
      adc_rom[3310] <= 8185;
      adc_rom[3311] <= 8186;
      adc_rom[3312] <= 8186;
      adc_rom[3313] <= 8188;
      adc_rom[3314] <= 8188;
      adc_rom[3315] <= 8187;
      adc_rom[3316] <= 8186;
      adc_rom[3317] <= 8186;
      adc_rom[3318] <= 8185;
      adc_rom[3319] <= 8188;
      adc_rom[3320] <= 8185;
      adc_rom[3321] <= 8187;
      adc_rom[3322] <= 8187;
      adc_rom[3323] <= 8187;
      adc_rom[3324] <= 8187;
      adc_rom[3325] <= 8186;
      adc_rom[3326] <= 8188;
      adc_rom[3327] <= 8189;
      adc_rom[3328] <= 8186;
      adc_rom[3329] <= 8188;
      adc_rom[3330] <= 8186;
      adc_rom[3331] <= 8187;
      adc_rom[3332] <= 8189;
      adc_rom[3333] <= 8184;
      adc_rom[3334] <= 8186;
      adc_rom[3335] <= 8184;
      adc_rom[3336] <= 8186;
      adc_rom[3337] <= 8186;
      adc_rom[3338] <= 8185;
      adc_rom[3339] <= 8187;
      adc_rom[3340] <= 8186;
      adc_rom[3341] <= 8185;
      adc_rom[3342] <= 8185;
      adc_rom[3343] <= 8187;
      adc_rom[3344] <= 8186;
      adc_rom[3345] <= 8187;
      adc_rom[3346] <= 8186;
      adc_rom[3347] <= 8187;
      adc_rom[3348] <= 8186;
      adc_rom[3349] <= 8187;
      adc_rom[3350] <= 8185;
      adc_rom[3351] <= 8186;
      adc_rom[3352] <= 8187;
      adc_rom[3353] <= 8185;
      adc_rom[3354] <= 8187;
      adc_rom[3355] <= 8186;
      adc_rom[3356] <= 8187;
      adc_rom[3357] <= 8188;
      adc_rom[3358] <= 8185;
      adc_rom[3359] <= 8188;
      adc_rom[3360] <= 8186;
      adc_rom[3361] <= 8187;
      adc_rom[3362] <= 8186;
      adc_rom[3363] <= 8185;
      adc_rom[3364] <= 8185;
      adc_rom[3365] <= 8186;
      adc_rom[3366] <= 8185;
      adc_rom[3367] <= 8185;
      adc_rom[3368] <= 8185;
      adc_rom[3369] <= 8186;
      adc_rom[3370] <= 8187;
      adc_rom[3371] <= 8185;
      adc_rom[3372] <= 8187;
      adc_rom[3373] <= 8185;
      adc_rom[3374] <= 8186;
      adc_rom[3375] <= 8185;
      adc_rom[3376] <= 8186;
      adc_rom[3377] <= 8186;
      adc_rom[3378] <= 8187;
      adc_rom[3379] <= 8186;
      adc_rom[3380] <= 8185;
      adc_rom[3381] <= 8186;
      adc_rom[3382] <= 8186;
      adc_rom[3383] <= 8185;
      adc_rom[3384] <= 8186;
      adc_rom[3385] <= 8186;
      adc_rom[3386] <= 8185;
      adc_rom[3387] <= 8185;
      adc_rom[3388] <= 8185;
      adc_rom[3389] <= 8189;
      adc_rom[3390] <= 8186;
      adc_rom[3391] <= 8186;
      adc_rom[3392] <= 8187;
      adc_rom[3393] <= 8185;
      adc_rom[3394] <= 8186;
      adc_rom[3395] <= 8186;
      adc_rom[3396] <= 8187;
      adc_rom[3397] <= 8187;
      adc_rom[3398] <= 8184;
      adc_rom[3399] <= 8187;
      adc_rom[3400] <= 8186;
      adc_rom[3401] <= 8188;
      adc_rom[3402] <= 8187;
      adc_rom[3403] <= 8187;
      adc_rom[3404] <= 8186;
      adc_rom[3405] <= 8188;
      adc_rom[3406] <= 8186;
      adc_rom[3407] <= 8188;
      adc_rom[3408] <= 8185;
      adc_rom[3409] <= 8187;
      adc_rom[3410] <= 8187;
      adc_rom[3411] <= 8187;
      adc_rom[3412] <= 8188;
      adc_rom[3413] <= 8184;
      adc_rom[3414] <= 8185;
      adc_rom[3415] <= 8184;
      adc_rom[3416] <= 8187;
      adc_rom[3417] <= 8187;
      adc_rom[3418] <= 8186;
      adc_rom[3419] <= 8187;
      adc_rom[3420] <= 8186;
      adc_rom[3421] <= 8188;
      adc_rom[3422] <= 8186;
      adc_rom[3423] <= 8185;
      adc_rom[3424] <= 8186;
      adc_rom[3425] <= 8186;
      adc_rom[3426] <= 8186;
      adc_rom[3427] <= 8187;
      adc_rom[3428] <= 8185;
      adc_rom[3429] <= 8187;
      adc_rom[3430] <= 8185;
      adc_rom[3431] <= 8186;
      adc_rom[3432] <= 8187;
      adc_rom[3433] <= 8184;
      adc_rom[3434] <= 8188;
      adc_rom[3435] <= 8186;
      adc_rom[3436] <= 8188;
      adc_rom[3437] <= 8187;
      adc_rom[3438] <= 8184;
      adc_rom[3439] <= 8188;
      adc_rom[3440] <= 8184;
      adc_rom[3441] <= 8188;
      adc_rom[3442] <= 8189;
      adc_rom[3443] <= 8186;
      adc_rom[3444] <= 8187;
      adc_rom[3445] <= 8188;
      adc_rom[3446] <= 8188;
      adc_rom[3447] <= 8187;
      adc_rom[3448] <= 8185;
      adc_rom[3449] <= 8187;
      adc_rom[3450] <= 8186;
      adc_rom[3451] <= 8188;
      adc_rom[3452] <= 8187;
      adc_rom[3453] <= 8186;
      adc_rom[3454] <= 8187;
      adc_rom[3455] <= 8185;
      adc_rom[3456] <= 8185;
      adc_rom[3457] <= 8187;
      adc_rom[3458] <= 8186;
      adc_rom[3459] <= 8188;
      adc_rom[3460] <= 8187;
      adc_rom[3461] <= 8188;
      adc_rom[3462] <= 8187;
      adc_rom[3463] <= 8187;
      adc_rom[3464] <= 8188;
      adc_rom[3465] <= 8186;
      adc_rom[3466] <= 8186;
      adc_rom[3467] <= 8188;
      adc_rom[3468] <= 8187;
      adc_rom[3469] <= 8188;
      adc_rom[3470] <= 8187;
      adc_rom[3471] <= 8187;
      adc_rom[3472] <= 8190;
      adc_rom[3473] <= 8186;
      adc_rom[3474] <= 8187;
      adc_rom[3475] <= 8187;
      adc_rom[3476] <= 8188;
      adc_rom[3477] <= 8187;
      adc_rom[3478] <= 8187;
      adc_rom[3479] <= 8188;
      adc_rom[3480] <= 8187;
      adc_rom[3481] <= 8187;
      adc_rom[3482] <= 8187;
      adc_rom[3483] <= 8186;
      adc_rom[3484] <= 8187;
      adc_rom[3485] <= 8187;
      adc_rom[3486] <= 8186;
      adc_rom[3487] <= 8187;
      adc_rom[3488] <= 8186;
      adc_rom[3489] <= 8187;
      adc_rom[3490] <= 8187;
      adc_rom[3491] <= 8187;
      adc_rom[3492] <= 8189;
      adc_rom[3493] <= 8185;
      adc_rom[3494] <= 8188;
      adc_rom[3495] <= 8187;
      adc_rom[3496] <= 8186;
      adc_rom[3497] <= 8188;
      adc_rom[3498] <= 8185;
      adc_rom[3499] <= 8188;
      adc_rom[3500] <= 8186;
      adc_rom[3501] <= 8185;
      adc_rom[3502] <= 8187;
      adc_rom[3503] <= 8186;
      adc_rom[3504] <= 8186;
      adc_rom[3505] <= 8185;
      adc_rom[3506] <= 8185;
      adc_rom[3507] <= 8189;
      adc_rom[3508] <= 8185;
      adc_rom[3509] <= 8188;
      adc_rom[3510] <= 8185;
      adc_rom[3511] <= 8186;
      adc_rom[3512] <= 8189;
      adc_rom[3513] <= 8186;
      adc_rom[3514] <= 8188;
      adc_rom[3515] <= 8186;
      adc_rom[3516] <= 8185;
      adc_rom[3517] <= 8188;
      adc_rom[3518] <= 8185;
      adc_rom[3519] <= 8188;
      adc_rom[3520] <= 8187;
      adc_rom[3521] <= 8187;
      adc_rom[3522] <= 8189;
      adc_rom[3523] <= 8186;
      adc_rom[3524] <= 8187;
      adc_rom[3525] <= 8185;
      adc_rom[3526] <= 8187;
      adc_rom[3527] <= 8188;
      adc_rom[3528] <= 8186;
      adc_rom[3529] <= 8185;
      adc_rom[3530] <= 8185;
      adc_rom[3531] <= 8188;
      adc_rom[3532] <= 8187;
      adc_rom[3533] <= 8187;
      adc_rom[3534] <= 8186;
      adc_rom[3535] <= 8186;
      adc_rom[3536] <= 8188;
      adc_rom[3537] <= 8188;
      adc_rom[3538] <= 8186;
      adc_rom[3539] <= 8188;
      adc_rom[3540] <= 8186;
      adc_rom[3541] <= 8187;
      adc_rom[3542] <= 8188;
      adc_rom[3543] <= 8185;
      adc_rom[3544] <= 8188;
      adc_rom[3545] <= 8187;
      adc_rom[3546] <= 8186;
      adc_rom[3547] <= 8187;
      adc_rom[3548] <= 8186;
      adc_rom[3549] <= 8187;
      adc_rom[3550] <= 8185;
      adc_rom[3551] <= 8189;
      adc_rom[3552] <= 8187;
      adc_rom[3553] <= 8186;
      adc_rom[3554] <= 8187;
      adc_rom[3555] <= 8186;
      adc_rom[3556] <= 8187;
      adc_rom[3557] <= 8185;
      adc_rom[3558] <= 8186;
      adc_rom[3559] <= 8188;
      adc_rom[3560] <= 8186;
      adc_rom[3561] <= 8185;
      adc_rom[3562] <= 8185;
      adc_rom[3563] <= 8185;
      adc_rom[3564] <= 8186;
      adc_rom[3565] <= 8186;
      adc_rom[3566] <= 8188;
      adc_rom[3567] <= 8187;
      adc_rom[3568] <= 8184;
      adc_rom[3569] <= 8187;
      adc_rom[3570] <= 8186;
      adc_rom[3571] <= 8184;
      adc_rom[3572] <= 8187;
      adc_rom[3573] <= 8186;
      adc_rom[3574] <= 8185;
      adc_rom[3575] <= 8185;
      adc_rom[3576] <= 8187;
      adc_rom[3577] <= 8188;
      adc_rom[3578] <= 8186;
      adc_rom[3579] <= 8187;
      adc_rom[3580] <= 8186;
      adc_rom[3581] <= 8184;
      adc_rom[3582] <= 8188;
      adc_rom[3583] <= 8186;
      adc_rom[3584] <= 8187;
      adc_rom[3585] <= 8187;
      adc_rom[3586] <= 8186;
      adc_rom[3587] <= 8187;
      adc_rom[3588] <= 8186;
      adc_rom[3589] <= 8187;
      adc_rom[3590] <= 8187;
      adc_rom[3591] <= 8187;
      adc_rom[3592] <= 8187;
      adc_rom[3593] <= 8186;
      adc_rom[3594] <= 8189;
      adc_rom[3595] <= 8186;
      adc_rom[3596] <= 8186;
      adc_rom[3597] <= 8184;
      adc_rom[3598] <= 8186;
      adc_rom[3599] <= 8188;
      adc_rom[3600] <= 8187;
      adc_rom[3601] <= 8186;
      adc_rom[3602] <= 8187;
      adc_rom[3603] <= 8186;
      adc_rom[3604] <= 8188;
      adc_rom[3605] <= 8186;
      adc_rom[3606] <= 8185;
      adc_rom[3607] <= 8186;
      adc_rom[3608] <= 8185;
      adc_rom[3609] <= 8187;
      adc_rom[3610] <= 8186;
      adc_rom[3611] <= 8186;
      adc_rom[3612] <= 8185;
      adc_rom[3613] <= 8186;
      adc_rom[3614] <= 8187;
      adc_rom[3615] <= 8185;
      adc_rom[3616] <= 8187;
      adc_rom[3617] <= 8189;
      adc_rom[3618] <= 8185;
      adc_rom[3619] <= 8186;
      adc_rom[3620] <= 8187;
      adc_rom[3621] <= 8187;
      adc_rom[3622] <= 8187;
      adc_rom[3623] <= 8185;
      adc_rom[3624] <= 8188;
      adc_rom[3625] <= 8186;
      adc_rom[3626] <= 8187;
      adc_rom[3627] <= 8188;
      adc_rom[3628] <= 8186;
      adc_rom[3629] <= 8186;
      adc_rom[3630] <= 8186;
      adc_rom[3631] <= 8187;
      adc_rom[3632] <= 8187;
      adc_rom[3633] <= 8185;
      adc_rom[3634] <= 8188;
      adc_rom[3635] <= 8188;
      adc_rom[3636] <= 8184;
      adc_rom[3637] <= 8188;
      adc_rom[3638] <= 8185;
      adc_rom[3639] <= 8187;
      adc_rom[3640] <= 8185;
      adc_rom[3641] <= 8185;
      adc_rom[3642] <= 8188;
      adc_rom[3643] <= 8184;
      adc_rom[3644] <= 8188;
      adc_rom[3645] <= 8186;
      adc_rom[3646] <= 8185;
      adc_rom[3647] <= 8189;
      adc_rom[3648] <= 8185;
      adc_rom[3649] <= 8187;
      adc_rom[3650] <= 8185;
      adc_rom[3651] <= 8187;
      adc_rom[3652] <= 8187;
      adc_rom[3653] <= 8187;
      adc_rom[3654] <= 8189;
      adc_rom[3655] <= 8185;
      adc_rom[3656] <= 8188;
      adc_rom[3657] <= 8185;
      adc_rom[3658] <= 8185;
      adc_rom[3659] <= 8187;
      adc_rom[3660] <= 8184;
      adc_rom[3661] <= 8187;
      adc_rom[3662] <= 8189;
      adc_rom[3663] <= 8187;
      adc_rom[3664] <= 8188;
      adc_rom[3665] <= 8187;
      adc_rom[3666] <= 8186;
      adc_rom[3667] <= 8190;
      adc_rom[3668] <= 8185;
      adc_rom[3669] <= 8187;
      adc_rom[3670] <= 8185;
      adc_rom[3671] <= 8187;
      adc_rom[3672] <= 8188;
      adc_rom[3673] <= 8187;
      adc_rom[3674] <= 8187;
      adc_rom[3675] <= 8185;
      adc_rom[3676] <= 8185;
      adc_rom[3677] <= 8187;
      adc_rom[3678] <= 8185;
      adc_rom[3679] <= 8187;
      adc_rom[3680] <= 8186;
      adc_rom[3681] <= 8187;
      adc_rom[3682] <= 8187;
      adc_rom[3683] <= 8187;
      adc_rom[3684] <= 8188;
      adc_rom[3685] <= 8189;
      adc_rom[3686] <= 8187;
      adc_rom[3687] <= 8187;
      adc_rom[3688] <= 8185;
      adc_rom[3689] <= 8188;
      adc_rom[3690] <= 8186;
      adc_rom[3691] <= 8187;
      adc_rom[3692] <= 8186;
      adc_rom[3693] <= 8186;
      adc_rom[3694] <= 8191;
      adc_rom[3695] <= 8187;
      adc_rom[3696] <= 8187;
      adc_rom[3697] <= 8186;
      adc_rom[3698] <= 8187;
      adc_rom[3699] <= 8186;
      adc_rom[3700] <= 8189;
      adc_rom[3701] <= 8188;
      adc_rom[3702] <= 8190;
      adc_rom[3703] <= 8186;
      adc_rom[3704] <= 8187;
      adc_rom[3705] <= 8187;
      adc_rom[3706] <= 8188;
      adc_rom[3707] <= 8189;
      adc_rom[3708] <= 8186;
      adc_rom[3709] <= 8187;
      adc_rom[3710] <= 8185;
      adc_rom[3711] <= 8188;
      adc_rom[3712] <= 8187;
      adc_rom[3713] <= 8187;
      adc_rom[3714] <= 8187;
      adc_rom[3715] <= 8184;
      adc_rom[3716] <= 8187;
      adc_rom[3717] <= 8187;
      adc_rom[3718] <= 8186;
      adc_rom[3719] <= 8188;
      adc_rom[3720] <= 8188;
      adc_rom[3721] <= 8187;
      adc_rom[3722] <= 8186;
      adc_rom[3723] <= 8187;
      adc_rom[3724] <= 8187;
      adc_rom[3725] <= 8186;
      adc_rom[3726] <= 8186;
      adc_rom[3727] <= 8187;
      adc_rom[3728] <= 8187;
      adc_rom[3729] <= 8188;
      adc_rom[3730] <= 8186;
      adc_rom[3731] <= 8187;
      adc_rom[3732] <= 8186;
      adc_rom[3733] <= 8185;
      adc_rom[3734] <= 8187;
      adc_rom[3735] <= 8185;
      adc_rom[3736] <= 8188;
      adc_rom[3737] <= 8186;
      adc_rom[3738] <= 8184;
      adc_rom[3739] <= 8186;
      adc_rom[3740] <= 8189;
      adc_rom[3741] <= 8188;
      adc_rom[3742] <= 8188;
      adc_rom[3743] <= 8186;
      adc_rom[3744] <= 8185;
      adc_rom[3745] <= 8186;
      adc_rom[3746] <= 8189;
      adc_rom[3747] <= 8189;
      adc_rom[3748] <= 8187;
      adc_rom[3749] <= 8187;
      adc_rom[3750] <= 8186;
      adc_rom[3751] <= 8187;
      adc_rom[3752] <= 8187;
      adc_rom[3753] <= 8186;
      adc_rom[3754] <= 8187;
      adc_rom[3755] <= 8186;
      adc_rom[3756] <= 8186;
      adc_rom[3757] <= 8185;
      adc_rom[3758] <= 8185;
      adc_rom[3759] <= 8189;
      adc_rom[3760] <= 8186;
      adc_rom[3761] <= 8187;
      adc_rom[3762] <= 8187;
      adc_rom[3763] <= 8185;
      adc_rom[3764] <= 8188;
      adc_rom[3765] <= 8187;
      adc_rom[3766] <= 8186;
      adc_rom[3767] <= 8189;
      adc_rom[3768] <= 8185;
      adc_rom[3769] <= 8187;
      adc_rom[3770] <= 8187;
      adc_rom[3771] <= 8187;
      adc_rom[3772] <= 8186;
      adc_rom[3773] <= 8186;
      adc_rom[3774] <= 8187;
      adc_rom[3775] <= 8185;
      adc_rom[3776] <= 8187;
      adc_rom[3777] <= 8187;
      adc_rom[3778] <= 8188;
      adc_rom[3779] <= 8188;
      adc_rom[3780] <= 8185;
      adc_rom[3781] <= 8185;
      adc_rom[3782] <= 8186;
      adc_rom[3783] <= 8187;
      adc_rom[3784] <= 8188;
      adc_rom[3785] <= 8185;
      adc_rom[3786] <= 8187;
      adc_rom[3787] <= 8185;
      adc_rom[3788] <= 8187;
      adc_rom[3789] <= 8187;
      adc_rom[3790] <= 8184;
      adc_rom[3791] <= 8186;
      adc_rom[3792] <= 8186;
      adc_rom[3793] <= 8185;
      adc_rom[3794] <= 8185;
      adc_rom[3795] <= 8185;
      adc_rom[3796] <= 8185;
      adc_rom[3797] <= 8186;
      adc_rom[3798] <= 8186;
      adc_rom[3799] <= 8186;
      adc_rom[3800] <= 8186;
      adc_rom[3801] <= 8186;
      adc_rom[3802] <= 8187;
      adc_rom[3803] <= 8187;
      adc_rom[3804] <= 8186;
      adc_rom[3805] <= 8187;
      adc_rom[3806] <= 8186;
      adc_rom[3807] <= 8187;
      adc_rom[3808] <= 8187;
      adc_rom[3809] <= 8188;
      adc_rom[3810] <= 8187;
      adc_rom[3811] <= 8187;
      adc_rom[3812] <= 8188;
      adc_rom[3813] <= 8188;
      adc_rom[3814] <= 8188;
      adc_rom[3815] <= 8187;
      adc_rom[3816] <= 8188;
      adc_rom[3817] <= 8188;
      adc_rom[3818] <= 8186;
      adc_rom[3819] <= 8188;
      adc_rom[3820] <= 8187;
      adc_rom[3821] <= 8188;
      adc_rom[3822] <= 8186;
      adc_rom[3823] <= 8187;
      adc_rom[3824] <= 8188;
      adc_rom[3825] <= 8185;
      adc_rom[3826] <= 8188;
      adc_rom[3827] <= 8189;
      adc_rom[3828] <= 8185;
      adc_rom[3829] <= 8187;
      adc_rom[3830] <= 8188;
      adc_rom[3831] <= 8188;
      adc_rom[3832] <= 8188;
      adc_rom[3833] <= 8185;
      adc_rom[3834] <= 8187;
      adc_rom[3835] <= 8185;
      adc_rom[3836] <= 8186;
      adc_rom[3837] <= 8187;
      adc_rom[3838] <= 8185;
      adc_rom[3839] <= 8190;
      adc_rom[3840] <= 8186;
      adc_rom[3841] <= 8187;
      adc_rom[3842] <= 8187;
      adc_rom[3843] <= 8186;
      adc_rom[3844] <= 8188;
      adc_rom[3845] <= 8186;
      adc_rom[3846] <= 8189;
      adc_rom[3847] <= 8189;
      adc_rom[3848] <= 8186;
      adc_rom[3849] <= 8187;
      adc_rom[3850] <= 8186;
      adc_rom[3851] <= 8190;
      adc_rom[3852] <= 8189;
      adc_rom[3853] <= 8185;
      adc_rom[3854] <= 8186;
      adc_rom[3855] <= 8184;
      adc_rom[3856] <= 8187;
      adc_rom[3857] <= 8187;
      adc_rom[3858] <= 8185;
      adc_rom[3859] <= 8187;
      adc_rom[3860] <= 8186;
      adc_rom[3861] <= 8187;
      adc_rom[3862] <= 8188;
      adc_rom[3863] <= 8187;
      adc_rom[3864] <= 8189;
      adc_rom[3865] <= 8188;
      adc_rom[3866] <= 8187;
      adc_rom[3867] <= 8187;
      adc_rom[3868] <= 8186;
      adc_rom[3869] <= 8189;
      adc_rom[3870] <= 8186;
      adc_rom[3871] <= 8186;
      adc_rom[3872] <= 8187;
      adc_rom[3873] <= 8187;
      adc_rom[3874] <= 8189;
      adc_rom[3875] <= 8186;
      adc_rom[3876] <= 8186;
      adc_rom[3877] <= 8190;
      adc_rom[3878] <= 8187;
      adc_rom[3879] <= 8187;
      adc_rom[3880] <= 8188;
      adc_rom[3881] <= 8188;
      adc_rom[3882] <= 8189;
      adc_rom[3883] <= 8185;
      adc_rom[3884] <= 8187;
      adc_rom[3885] <= 8187;
      adc_rom[3886] <= 8184;
      adc_rom[3887] <= 8186;
      adc_rom[3888] <= 8184;
      adc_rom[3889] <= 8187;
      adc_rom[3890] <= 8187;
      adc_rom[3891] <= 8185;
      adc_rom[3892] <= 8186;
      adc_rom[3893] <= 8185;
      adc_rom[3894] <= 8188;
      adc_rom[3895] <= 8186;
      adc_rom[3896] <= 8187;
      adc_rom[3897] <= 8188;
      adc_rom[3898] <= 8188;
      adc_rom[3899] <= 8187;
      adc_rom[3900] <= 8186;
      adc_rom[3901] <= 8187;
      adc_rom[3902] <= 8186;
      adc_rom[3903] <= 8186;
      adc_rom[3904] <= 8187;
      adc_rom[3905] <= 8185;
      adc_rom[3906] <= 8188;
      adc_rom[3907] <= 8187;
      adc_rom[3908] <= 8184;
      adc_rom[3909] <= 8186;
      adc_rom[3910] <= 8187;
      adc_rom[3911] <= 8188;
      adc_rom[3912] <= 8189;
      adc_rom[3913] <= 8187;
      adc_rom[3914] <= 8187;
      adc_rom[3915] <= 8186;
      adc_rom[3916] <= 8186;
      adc_rom[3917] <= 8187;
      adc_rom[3918] <= 8186;
      adc_rom[3919] <= 8187;
      adc_rom[3920] <= 8186;
      adc_rom[3921] <= 8188;
      adc_rom[3922] <= 8189;
      adc_rom[3923] <= 8186;
      adc_rom[3924] <= 8189;
      adc_rom[3925] <= 8186;
      adc_rom[3926] <= 8187;
      adc_rom[3927] <= 8186;
      adc_rom[3928] <= 8186;
      adc_rom[3929] <= 8187;
      adc_rom[3930] <= 8187;
      adc_rom[3931] <= 8187;
      adc_rom[3932] <= 8186;
      adc_rom[3933] <= 8188;
      adc_rom[3934] <= 8188;
      adc_rom[3935] <= 8187;
      adc_rom[3936] <= 8189;
      adc_rom[3937] <= 8186;
      adc_rom[3938] <= 8188;
      adc_rom[3939] <= 8189;
      adc_rom[3940] <= 8186;
      adc_rom[3941] <= 8188;
      adc_rom[3942] <= 8189;
      adc_rom[3943] <= 8187;
      adc_rom[3944] <= 8187;
      adc_rom[3945] <= 8185;
      adc_rom[3946] <= 8187;
      adc_rom[3947] <= 8187;
      adc_rom[3948] <= 8185;
      adc_rom[3949] <= 8189;
      adc_rom[3950] <= 8186;
      adc_rom[3951] <= 8187;
      adc_rom[3952] <= 8188;
      adc_rom[3953] <= 8188;
      adc_rom[3954] <= 8187;
      adc_rom[3955] <= 8186;
      adc_rom[3956] <= 8189;
      adc_rom[3957] <= 8187;
      adc_rom[3958] <= 8186;
      adc_rom[3959] <= 8189;
      adc_rom[3960] <= 8189;
      adc_rom[3961] <= 8187;
      adc_rom[3962] <= 8189;
      adc_rom[3963] <= 8185;
      adc_rom[3964] <= 8188;
      adc_rom[3965] <= 8186;
      adc_rom[3966] <= 8188;
      adc_rom[3967] <= 8187;
      adc_rom[3968] <= 8184;
      adc_rom[3969] <= 8188;
      adc_rom[3970] <= 8186;
      adc_rom[3971] <= 8187;
      adc_rom[3972] <= 8187;
      adc_rom[3973] <= 8188;
      adc_rom[3974] <= 8187;
      adc_rom[3975] <= 8184;
      adc_rom[3976] <= 8186;
      adc_rom[3977] <= 8187;
      adc_rom[3978] <= 8187;
      adc_rom[3979] <= 8187;
      adc_rom[3980] <= 8185;
      adc_rom[3981] <= 8186;
      adc_rom[3982] <= 8188;
      adc_rom[3983] <= 8187;
      adc_rom[3984] <= 8186;
      adc_rom[3985] <= 8186;
      adc_rom[3986] <= 8189;
      adc_rom[3987] <= 8188;
      adc_rom[3988] <= 8185;
      adc_rom[3989] <= 8187;
      adc_rom[3990] <= 8186;
      adc_rom[3991] <= 8187;
      adc_rom[3992] <= 8188;
      adc_rom[3993] <= 8185;
      adc_rom[3994] <= 8187;
      adc_rom[3995] <= 8187;
      adc_rom[3996] <= 8187;
      adc_rom[3997] <= 8187;
      adc_rom[3998] <= 8187;
      adc_rom[3999] <= 8187;
      adc_rom[4000] <= 8189;
      adc_rom[4001] <= 8186;
      adc_rom[4002] <= 8187;
      adc_rom[4003] <= 8187;
      adc_rom[4004] <= 8188;
      adc_rom[4005] <= 8186;
      adc_rom[4006] <= 8186;
      adc_rom[4007] <= 8188;
      adc_rom[4008] <= 8186;
      adc_rom[4009] <= 8189;
      adc_rom[4010] <= 8187;
      adc_rom[4011] <= 8187;
      adc_rom[4012] <= 8186;
      adc_rom[4013] <= 8186;
      adc_rom[4014] <= 8186;
      adc_rom[4015] <= 8186;
      adc_rom[4016] <= 8186;
      adc_rom[4017] <= 8188;
      adc_rom[4018] <= 8187;
      adc_rom[4019] <= 8189;
      adc_rom[4020] <= 8186;
      adc_rom[4021] <= 8186;
      adc_rom[4022] <= 8189;
      adc_rom[4023] <= 8188;
      adc_rom[4024] <= 8189;
      adc_rom[4025] <= 8184;
      adc_rom[4026] <= 8190;
      adc_rom[4027] <= 8187;
      adc_rom[4028] <= 8188;
      adc_rom[4029] <= 8187;
      adc_rom[4030] <= 8185;
      adc_rom[4031] <= 8187;
      adc_rom[4032] <= 8189;
      adc_rom[4033] <= 8186;
      adc_rom[4034] <= 8187;
      adc_rom[4035] <= 8185;
      adc_rom[4036] <= 8187;
      adc_rom[4037] <= 8187;
      adc_rom[4038] <= 8187;
      adc_rom[4039] <= 8188;
      adc_rom[4040] <= 8187;
      adc_rom[4041] <= 8186;
      adc_rom[4042] <= 8189;
      adc_rom[4043] <= 8186;
      adc_rom[4044] <= 8189;
      adc_rom[4045] <= 8189;
      adc_rom[4046] <= 8187;
      adc_rom[4047] <= 8189;
      adc_rom[4048] <= 8188;
      adc_rom[4049] <= 8185;
      adc_rom[4050] <= 8186;
      adc_rom[4051] <= 8188;
      adc_rom[4052] <= 8188;
      adc_rom[4053] <= 8187;
      adc_rom[4054] <= 8187;
      adc_rom[4055] <= 8187;
      adc_rom[4056] <= 8186;
      adc_rom[4057] <= 8189;
      adc_rom[4058] <= 8188;
      adc_rom[4059] <= 8188;
      adc_rom[4060] <= 8185;
      adc_rom[4061] <= 8188;
      adc_rom[4062] <= 8187;
      adc_rom[4063] <= 8185;
      adc_rom[4064] <= 8187;
      adc_rom[4065] <= 8187;
      adc_rom[4066] <= 8187;
      adc_rom[4067] <= 8189;
      adc_rom[4068] <= 8185;
      adc_rom[4069] <= 8187;
      adc_rom[4070] <= 8184;
      adc_rom[4071] <= 8185;
      adc_rom[4072] <= 8188;
      adc_rom[4073] <= 8185;
      adc_rom[4074] <= 8186;
      adc_rom[4075] <= 8185;
      adc_rom[4076] <= 8187;
      adc_rom[4077] <= 8188;
      adc_rom[4078] <= 8188;
      adc_rom[4079] <= 8187;
      adc_rom[4080] <= 8185;
      adc_rom[4081] <= 8187;
      adc_rom[4082] <= 8187;
      adc_rom[4083] <= 8186;
      adc_rom[4084] <= 8186;
      adc_rom[4085] <= 8188;
      adc_rom[4086] <= 8185;
      adc_rom[4087] <= 8187;
      adc_rom[4088] <= 8189;
      adc_rom[4089] <= 8185;
      adc_rom[4090] <= 8187;
      adc_rom[4091] <= 8187;
      adc_rom[4092] <= 8184;
      adc_rom[4093] <= 8188;
      adc_rom[4094] <= 8187;
      adc_rom[4095] <= 8185;
      adc_rom[4096] <= 8190;
      adc_rom[4097] <= 8186;
      adc_rom[4098] <= 8186;
      adc_rom[4099] <= 8187;
      adc_rom[4100] <= 8186;
      adc_rom[4101] <= 8188;
      adc_rom[4102] <= 8187;
      adc_rom[4103] <= 8187;
      adc_rom[4104] <= 8189;
      adc_rom[4105] <= 8186;
      adc_rom[4106] <= 8187;
      adc_rom[4107] <= 8185;
      adc_rom[4108] <= 8185;
      adc_rom[4109] <= 8187;
      adc_rom[4110] <= 8187;
      adc_rom[4111] <= 8187;
      adc_rom[4112] <= 8188;
      adc_rom[4113] <= 8186;
      adc_rom[4114] <= 8186;
      adc_rom[4115] <= 8185;
      adc_rom[4116] <= 8187;
      adc_rom[4117] <= 8187;
      adc_rom[4118] <= 8183;
      adc_rom[4119] <= 8187;
      adc_rom[4120] <= 8183;
      adc_rom[4121] <= 8186;
      adc_rom[4122] <= 8186;
      adc_rom[4123] <= 8184;
      adc_rom[4124] <= 8188;
      adc_rom[4125] <= 8186;
      adc_rom[4126] <= 8185;
      adc_rom[4127] <= 8187;
      adc_rom[4128] <= 8185;
      adc_rom[4129] <= 8189;
      adc_rom[4130] <= 8187;
      adc_rom[4131] <= 8187;
      adc_rom[4132] <= 8187;
      adc_rom[4133] <= 8187;
      adc_rom[4134] <= 8188;
      adc_rom[4135] <= 8187;
      adc_rom[4136] <= 8187;
      adc_rom[4137] <= 8186;
      adc_rom[4138] <= 8187;
      adc_rom[4139] <= 8186;
      adc_rom[4140] <= 8186;
      adc_rom[4141] <= 8186;
      adc_rom[4142] <= 8187;
      adc_rom[4143] <= 8187;
      adc_rom[4144] <= 8187;
      adc_rom[4145] <= 8186;
      adc_rom[4146] <= 8186;
      adc_rom[4147] <= 8186;
      adc_rom[4148] <= 8187;
      adc_rom[4149] <= 8187;
      adc_rom[4150] <= 8185;
      adc_rom[4151] <= 8185;
      adc_rom[4152] <= 8188;
      adc_rom[4153] <= 8188;
      adc_rom[4154] <= 8188;
      adc_rom[4155] <= 8185;
      adc_rom[4156] <= 8187;
      adc_rom[4157] <= 8187;
      adc_rom[4158] <= 8185;
      adc_rom[4159] <= 8186;
      adc_rom[4160] <= 8185;
      adc_rom[4161] <= 8189;
      adc_rom[4162] <= 8187;
      adc_rom[4163] <= 8185;
      adc_rom[4164] <= 8189;
      adc_rom[4165] <= 8186;
      adc_rom[4166] <= 8186;
      adc_rom[4167] <= 8187;
      adc_rom[4168] <= 8187;
      adc_rom[4169] <= 8186;
      adc_rom[4170] <= 8186;
      adc_rom[4171] <= 8188;
      adc_rom[4172] <= 8187;
      adc_rom[4173] <= 8186;
      adc_rom[4174] <= 8187;
      adc_rom[4175] <= 8188;
      adc_rom[4176] <= 8186;
      adc_rom[4177] <= 8188;
      adc_rom[4178] <= 8186;
      adc_rom[4179] <= 8189;
      adc_rom[4180] <= 8186;
      adc_rom[4181] <= 8185;
      adc_rom[4182] <= 8185;
      adc_rom[4183] <= 8186;
      adc_rom[4184] <= 8187;
      adc_rom[4185] <= 8185;
      adc_rom[4186] <= 8186;
      adc_rom[4187] <= 8186;
      adc_rom[4188] <= 8185;
      adc_rom[4189] <= 8187;
      adc_rom[4190] <= 8188;
      adc_rom[4191] <= 8187;
      adc_rom[4192] <= 8187;
      adc_rom[4193] <= 8185;
      adc_rom[4194] <= 8187;
      adc_rom[4195] <= 8184;
      adc_rom[4196] <= 8187;
      adc_rom[4197] <= 8189;
      adc_rom[4198] <= 8185;
      adc_rom[4199] <= 8187;
      adc_rom[4200] <= 8185;
      adc_rom[4201] <= 8189;
      adc_rom[4202] <= 8188;
      adc_rom[4203] <= 8185;
      adc_rom[4204] <= 8188;
      adc_rom[4205] <= 8186;
      adc_rom[4206] <= 8186;
      adc_rom[4207] <= 8187;
      adc_rom[4208] <= 8186;
      adc_rom[4209] <= 8189;
      adc_rom[4210] <= 8187;
      adc_rom[4211] <= 8187;
      adc_rom[4212] <= 8187;
      adc_rom[4213] <= 8186;
      adc_rom[4214] <= 8189;
      adc_rom[4215] <= 8186;
      adc_rom[4216] <= 8186;
      adc_rom[4217] <= 8184;
      adc_rom[4218] <= 8185;
      adc_rom[4219] <= 8187;
      adc_rom[4220] <= 8186;
      adc_rom[4221] <= 8186;
      adc_rom[4222] <= 8189;
      adc_rom[4223] <= 8186;
      adc_rom[4224] <= 8186;
      adc_rom[4225] <= 8187;
      adc_rom[4226] <= 8188;
      adc_rom[4227] <= 8187;
      adc_rom[4228] <= 8185;
      adc_rom[4229] <= 8187;
      adc_rom[4230] <= 8183;
      adc_rom[4231] <= 8187;
      adc_rom[4232] <= 8186;
      adc_rom[4233] <= 8186;
      adc_rom[4234] <= 8187;
      adc_rom[4235] <= 8187;
      adc_rom[4236] <= 8187;
      adc_rom[4237] <= 8189;
      adc_rom[4238] <= 8186;
      adc_rom[4239] <= 8187;
      adc_rom[4240] <= 8186;
      adc_rom[4241] <= 8186;
      adc_rom[4242] <= 8189;
      adc_rom[4243] <= 8186;
      adc_rom[4244] <= 8190;
      adc_rom[4245] <= 8186;
      adc_rom[4246] <= 8186;
      adc_rom[4247] <= 8190;
      adc_rom[4248] <= 8186;
      adc_rom[4249] <= 8188;
      adc_rom[4250] <= 8187;
      adc_rom[4251] <= 8186;
      adc_rom[4252] <= 8189;
      adc_rom[4253] <= 8186;
      adc_rom[4254] <= 8186;
      adc_rom[4255] <= 8185;
      adc_rom[4256] <= 8187;
      adc_rom[4257] <= 8186;
      adc_rom[4258] <= 8186;
      adc_rom[4259] <= 8187;
      adc_rom[4260] <= 8185;
      adc_rom[4261] <= 8186;
      adc_rom[4262] <= 8186;
      adc_rom[4263] <= 8186;
      adc_rom[4264] <= 8188;
      adc_rom[4265] <= 8186;
      adc_rom[4266] <= 8188;
      adc_rom[4267] <= 8186;
      adc_rom[4268] <= 8184;
      adc_rom[4269] <= 8188;
      adc_rom[4270] <= 8187;
      adc_rom[4271] <= 8189;
      adc_rom[4272] <= 8188;
      adc_rom[4273] <= 8187;
      adc_rom[4274] <= 8189;
      adc_rom[4275] <= 8188;
      adc_rom[4276] <= 8185;
      adc_rom[4277] <= 8186;
      adc_rom[4278] <= 8187;
      adc_rom[4279] <= 8192;
      adc_rom[4280] <= 8186;
      adc_rom[4281] <= 8188;
      adc_rom[4282] <= 8189;
      adc_rom[4283] <= 8186;
      adc_rom[4284] <= 8187;
      adc_rom[4285] <= 8187;
      adc_rom[4286] <= 8187;
      adc_rom[4287] <= 8188;
      adc_rom[4288] <= 8188;
      adc_rom[4289] <= 8190;
      adc_rom[4290] <= 8186;
      adc_rom[4291] <= 8186;
      adc_rom[4292] <= 8187;
      adc_rom[4293] <= 8185;
      adc_rom[4294] <= 8187;
      adc_rom[4295] <= 8186;
      adc_rom[4296] <= 8187;
      adc_rom[4297] <= 8187;
      adc_rom[4298] <= 8185;
      adc_rom[4299] <= 8187;
      adc_rom[4300] <= 8186;
      adc_rom[4301] <= 8187;
      adc_rom[4302] <= 8187;
      adc_rom[4303] <= 8186;
      adc_rom[4304] <= 8187;
      adc_rom[4305] <= 8186;
      adc_rom[4306] <= 8186;
      adc_rom[4307] <= 8186;
      adc_rom[4308] <= 8187;
      adc_rom[4309] <= 8188;
      adc_rom[4310] <= 8185;
      adc_rom[4311] <= 8187;
      adc_rom[4312] <= 8187;
      adc_rom[4313] <= 8187;
      adc_rom[4314] <= 8187;
      adc_rom[4315] <= 8185;
      adc_rom[4316] <= 8188;
      adc_rom[4317] <= 8187;
      adc_rom[4318] <= 8186;
      adc_rom[4319] <= 8186;
      adc_rom[4320] <= 8185;
      adc_rom[4321] <= 8187;
      adc_rom[4322] <= 8186;
      adc_rom[4323] <= 8185;
      adc_rom[4324] <= 8189;
      adc_rom[4325] <= 8186;
      adc_rom[4326] <= 8186;
      adc_rom[4327] <= 8188;
      adc_rom[4328] <= 8185;
      adc_rom[4329] <= 8189;
      adc_rom[4330] <= 8187;
      adc_rom[4331] <= 8187;
      adc_rom[4332] <= 8186;
      adc_rom[4333] <= 8187;
      adc_rom[4334] <= 8189;
      adc_rom[4335] <= 8186;
      adc_rom[4336] <= 8188;
      adc_rom[4337] <= 8187;
      adc_rom[4338] <= 8188;
      adc_rom[4339] <= 8187;
      adc_rom[4340] <= 8185;
      adc_rom[4341] <= 8186;
      adc_rom[4342] <= 8188;
      adc_rom[4343] <= 8185;
      adc_rom[4344] <= 8189;
      adc_rom[4345] <= 8186;
      adc_rom[4346] <= 8188;
      adc_rom[4347] <= 8188;
      adc_rom[4348] <= 8187;
      adc_rom[4349] <= 8185;
      adc_rom[4350] <= 8187;
      adc_rom[4351] <= 8187;
      adc_rom[4352] <= 8187;
      adc_rom[4353] <= 8185;
      adc_rom[4354] <= 8187;
      adc_rom[4355] <= 8186;
      adc_rom[4356] <= 8187;
      adc_rom[4357] <= 8186;
      adc_rom[4358] <= 8184;
      adc_rom[4359] <= 8187;
      adc_rom[4360] <= 8188;
      adc_rom[4361] <= 8186;
      adc_rom[4362] <= 8187;
      adc_rom[4363] <= 8185;
      adc_rom[4364] <= 8188;
      adc_rom[4365] <= 8186;
      adc_rom[4366] <= 8187;
      adc_rom[4367] <= 8189;
      adc_rom[4368] <= 8184;
      adc_rom[4369] <= 8185;
      adc_rom[4370] <= 8187;
      adc_rom[4371] <= 8187;
      adc_rom[4372] <= 8187;
      adc_rom[4373] <= 8185;
      adc_rom[4374] <= 8187;
      adc_rom[4375] <= 8185;
      adc_rom[4376] <= 8187;
      adc_rom[4377] <= 8186;
      adc_rom[4378] <= 8185;
      adc_rom[4379] <= 8187;
      adc_rom[4380] <= 8186;
      adc_rom[4381] <= 8187;
      adc_rom[4382] <= 8189;
      adc_rom[4383] <= 8185;
      adc_rom[4384] <= 8187;
      adc_rom[4385] <= 8185;
      adc_rom[4386] <= 8186;
      adc_rom[4387] <= 8187;
      adc_rom[4388] <= 8185;
      adc_rom[4389] <= 8187;
      adc_rom[4390] <= 8186;
      adc_rom[4391] <= 8186;
      adc_rom[4392] <= 8186;
      adc_rom[4393] <= 8184;
      adc_rom[4394] <= 8185;
      adc_rom[4395] <= 8185;
      adc_rom[4396] <= 8186;
      adc_rom[4397] <= 8187;
      adc_rom[4398] <= 8184;
      adc_rom[4399] <= 8185;
      adc_rom[4400] <= 8184;
      adc_rom[4401] <= 8186;
      adc_rom[4402] <= 8186;
      adc_rom[4403] <= 8183;
      adc_rom[4404] <= 8185;
      adc_rom[4405] <= 8185;
      adc_rom[4406] <= 8187;
      adc_rom[4407] <= 8188;
      adc_rom[4408] <= 8187;
      adc_rom[4409] <= 8188;
      adc_rom[4410] <= 8184;
      adc_rom[4411] <= 8187;
      adc_rom[4412] <= 8187;
      adc_rom[4413] <= 8185;
      adc_rom[4414] <= 8187;
      adc_rom[4415] <= 8187;
      adc_rom[4416] <= 8187;
      adc_rom[4417] <= 8184;
      adc_rom[4418] <= 8185;
      adc_rom[4419] <= 8188;
      adc_rom[4420] <= 8187;
      adc_rom[4421] <= 8186;
      adc_rom[4422] <= 8186;
      adc_rom[4423] <= 8184;
      adc_rom[4424] <= 8186;
      adc_rom[4425] <= 8184;
      adc_rom[4426] <= 8186;
      adc_rom[4427] <= 8187;
      adc_rom[4428] <= 8186;
      adc_rom[4429] <= 8187;
      adc_rom[4430] <= 8186;
      adc_rom[4431] <= 8185;
      adc_rom[4432] <= 8185;
      adc_rom[4433] <= 8185;
      adc_rom[4434] <= 8187;
      adc_rom[4435] <= 8183;
      adc_rom[4436] <= 8185;
      adc_rom[4437] <= 8188;
      adc_rom[4438] <= 8186;
      adc_rom[4439] <= 8188;
      adc_rom[4440] <= 8186;
      adc_rom[4441] <= 8187;
      adc_rom[4442] <= 8187;
      adc_rom[4443] <= 8186;
      adc_rom[4444] <= 8188;
      adc_rom[4445] <= 8185;
      adc_rom[4446] <= 8186;
      adc_rom[4447] <= 8186;
      adc_rom[4448] <= 8186;
      adc_rom[4449] <= 8188;
      adc_rom[4450] <= 8186;
      adc_rom[4451] <= 8188;
      adc_rom[4452] <= 8187;
      adc_rom[4453] <= 8187;
      adc_rom[4454] <= 8185;
      adc_rom[4455] <= 8184;
      adc_rom[4456] <= 8186;
      adc_rom[4457] <= 8186;
      adc_rom[4458] <= 8185;
      adc_rom[4459] <= 8187;
      adc_rom[4460] <= 8184;
      adc_rom[4461] <= 8186;
      adc_rom[4462] <= 8187;
      adc_rom[4463] <= 8185;
      adc_rom[4464] <= 8187;
      adc_rom[4465] <= 8189;
      adc_rom[4466] <= 8187;
      adc_rom[4467] <= 8185;
      adc_rom[4468] <= 8185;
      adc_rom[4469] <= 8186;
      adc_rom[4470] <= 8186;
      adc_rom[4471] <= 8185;
      adc_rom[4472] <= 8187;
      adc_rom[4473] <= 8185;
      adc_rom[4474] <= 8188;
      adc_rom[4475] <= 8187;
      adc_rom[4476] <= 8185;
      adc_rom[4477] <= 8186;
      adc_rom[4478] <= 8187;
      adc_rom[4479] <= 8187;
      adc_rom[4480] <= 8186;
      adc_rom[4481] <= 8188;
      adc_rom[4482] <= 8188;
      adc_rom[4483] <= 8187;
      adc_rom[4484] <= 8188;
      adc_rom[4485] <= 8188;
      adc_rom[4486] <= 8186;
      adc_rom[4487] <= 8185;
      adc_rom[4488] <= 8185;
      adc_rom[4489] <= 8187;
      adc_rom[4490] <= 8186;
      adc_rom[4491] <= 8186;
      adc_rom[4492] <= 8189;
      adc_rom[4493] <= 8185;
      adc_rom[4494] <= 8188;
      adc_rom[4495] <= 8187;
      adc_rom[4496] <= 8187;
      adc_rom[4497] <= 8187;
      adc_rom[4498] <= 8185;
      adc_rom[4499] <= 8188;
      adc_rom[4500] <= 8185;
      adc_rom[4501] <= 8186;
      adc_rom[4502] <= 8189;
      adc_rom[4503] <= 8186;
      adc_rom[4504] <= 8187;
      adc_rom[4505] <= 8187;
      adc_rom[4506] <= 8187;
      adc_rom[4507] <= 8187;
      adc_rom[4508] <= 8186;
      adc_rom[4509] <= 8187;
      adc_rom[4510] <= 8186;
      adc_rom[4511] <= 8187;
      adc_rom[4512] <= 8189;
      adc_rom[4513] <= 8185;
      adc_rom[4514] <= 8187;
      adc_rom[4515] <= 8185;
      adc_rom[4516] <= 8187;
      adc_rom[4517] <= 8188;
      adc_rom[4518] <= 8186;
      adc_rom[4519] <= 8186;
      adc_rom[4520] <= 8187;
      adc_rom[4521] <= 8187;
      adc_rom[4522] <= 8186;
      adc_rom[4523] <= 8186;
      adc_rom[4524] <= 8188;
      adc_rom[4525] <= 8186;
      adc_rom[4526] <= 8186;
      adc_rom[4527] <= 8188;
      adc_rom[4528] <= 8185;
      adc_rom[4529] <= 8187;
      adc_rom[4530] <= 8186;
      adc_rom[4531] <= 8186;
      adc_rom[4532] <= 8188;
      adc_rom[4533] <= 8188;
      adc_rom[4534] <= 8187;
      adc_rom[4535] <= 8188;
      adc_rom[4536] <= 8186;
      adc_rom[4537] <= 8187;
      adc_rom[4538] <= 8187;
      adc_rom[4539] <= 8188;
      adc_rom[4540] <= 8185;
      adc_rom[4541] <= 8186;
      adc_rom[4542] <= 8187;
      adc_rom[4543] <= 8186;
      adc_rom[4544] <= 8188;
      adc_rom[4545] <= 8187;
      adc_rom[4546] <= 8188;
      adc_rom[4547] <= 8186;
      adc_rom[4548] <= 8184;
      adc_rom[4549] <= 8186;
      adc_rom[4550] <= 8185;
      adc_rom[4551] <= 8186;
      adc_rom[4552] <= 8189;
      adc_rom[4553] <= 8189;
      adc_rom[4554] <= 8189;
      adc_rom[4555] <= 8185;
      adc_rom[4556] <= 8186;
      adc_rom[4557] <= 8187;
      adc_rom[4558] <= 8185;
      adc_rom[4559] <= 8187;
      adc_rom[4560] <= 8185;
      adc_rom[4561] <= 8188;
      adc_rom[4562] <= 8187;
      adc_rom[4563] <= 8187;
      adc_rom[4564] <= 8189;
      adc_rom[4565] <= 8188;
      adc_rom[4566] <= 8188;
      adc_rom[4567] <= 8189;
      adc_rom[4568] <= 8187;
      adc_rom[4569] <= 8189;
      adc_rom[4570] <= 8186;
      adc_rom[4571] <= 8184;
      adc_rom[4572] <= 8188;
      adc_rom[4573] <= 8186;
      adc_rom[4574] <= 8188;
      adc_rom[4575] <= 8186;
      adc_rom[4576] <= 8186;
      adc_rom[4577] <= 8188;
      adc_rom[4578] <= 8186;
      adc_rom[4579] <= 8188;
      adc_rom[4580] <= 8186;
      adc_rom[4581] <= 8186;
      adc_rom[4582] <= 8187;
      adc_rom[4583] <= 8186;
      adc_rom[4584] <= 8187;
      adc_rom[4585] <= 8186;
      adc_rom[4586] <= 8189;
      adc_rom[4587] <= 8187;
      adc_rom[4588] <= 8186;
      adc_rom[4589] <= 8187;
      adc_rom[4590] <= 8187;
      adc_rom[4591] <= 8187;
      adc_rom[4592] <= 8186;
      adc_rom[4593] <= 8184;
      adc_rom[4594] <= 8187;
      adc_rom[4595] <= 8186;
      adc_rom[4596] <= 8186;
      adc_rom[4597] <= 8187;
      adc_rom[4598] <= 8185;
      adc_rom[4599] <= 8186;
      adc_rom[4600] <= 8187;
      adc_rom[4601] <= 8186;
      adc_rom[4602] <= 8187;
      adc_rom[4603] <= 8185;
      adc_rom[4604] <= 8188;
      adc_rom[4605] <= 8186;
      adc_rom[4606] <= 8186;
      adc_rom[4607] <= 8186;
      adc_rom[4608] <= 8187;
      adc_rom[4609] <= 8187;
      adc_rom[4610] <= 8187;
      adc_rom[4611] <= 8188;
      adc_rom[4612] <= 8188;
      adc_rom[4613] <= 8186;
      adc_rom[4614] <= 8187;
      adc_rom[4615] <= 8186;
      adc_rom[4616] <= 8186;
      adc_rom[4617] <= 8186;
      adc_rom[4618] <= 8186;
      adc_rom[4619] <= 8187;
      adc_rom[4620] <= 8186;
      adc_rom[4621] <= 8187;
      adc_rom[4622] <= 8187;
      adc_rom[4623] <= 8186;
      adc_rom[4624] <= 8186;
      adc_rom[4625] <= 8186;
      adc_rom[4626] <= 8186;
      adc_rom[4627] <= 8187;
      adc_rom[4628] <= 8185;
      adc_rom[4629] <= 8187;
      adc_rom[4630] <= 8186;
      adc_rom[4631] <= 8185;
      adc_rom[4632] <= 8189;
      adc_rom[4633] <= 8186;
      adc_rom[4634] <= 8189;
      adc_rom[4635] <= 8186;
      adc_rom[4636] <= 8187;
      adc_rom[4637] <= 8186;
      adc_rom[4638] <= 8185;
      adc_rom[4639] <= 8185;
      adc_rom[4640] <= 8186;
      adc_rom[4641] <= 8188;
      adc_rom[4642] <= 8188;
      adc_rom[4643] <= 8186;
      adc_rom[4644] <= 8187;
      adc_rom[4645] <= 8187;
      adc_rom[4646] <= 8188;
      adc_rom[4647] <= 8189;
      adc_rom[4648] <= 8186;
      adc_rom[4649] <= 8187;
      adc_rom[4650] <= 8186;
      adc_rom[4651] <= 8187;
      adc_rom[4652] <= 8188;
      adc_rom[4653] <= 8185;
      adc_rom[4654] <= 8188;
      adc_rom[4655] <= 8188;
      adc_rom[4656] <= 8189;
      adc_rom[4657] <= 8188;
      adc_rom[4658] <= 8188;
      adc_rom[4659] <= 8188;
      adc_rom[4660] <= 8186;
      adc_rom[4661] <= 8186;
      adc_rom[4662] <= 8187;
      adc_rom[4663] <= 8186;
      adc_rom[4664] <= 8188;
      adc_rom[4665] <= 8185;
      adc_rom[4666] <= 8188;
      adc_rom[4667] <= 8187;
      adc_rom[4668] <= 8185;
      adc_rom[4669] <= 8186;
      adc_rom[4670] <= 8187;
      adc_rom[4671] <= 8187;
      adc_rom[4672] <= 8188;
      adc_rom[4673] <= 8185;
      adc_rom[4674] <= 8185;
      adc_rom[4675] <= 8186;
      adc_rom[4676] <= 8187;
      adc_rom[4677] <= 8189;
      adc_rom[4678] <= 8187;
      adc_rom[4679] <= 8189;
      adc_rom[4680] <= 8185;
      adc_rom[4681] <= 8185;
      adc_rom[4682] <= 8187;
      adc_rom[4683] <= 8186;
      adc_rom[4684] <= 8187;
      adc_rom[4685] <= 8185;
      adc_rom[4686] <= 8188;
      adc_rom[4687] <= 8189;
      adc_rom[4688] <= 8186;
      adc_rom[4689] <= 8189;
      adc_rom[4690] <= 8186;
      adc_rom[4691] <= 8186;
      adc_rom[4692] <= 8188;
      adc_rom[4693] <= 8185;
      adc_rom[4694] <= 8187;
      adc_rom[4695] <= 8187;
      adc_rom[4696] <= 8187;
      adc_rom[4697] <= 8187;
      adc_rom[4698] <= 8185;
      adc_rom[4699] <= 8187;
      adc_rom[4700] <= 8186;
      adc_rom[4701] <= 8185;
      adc_rom[4702] <= 8187;
      adc_rom[4703] <= 8186;
      adc_rom[4704] <= 8185;
      adc_rom[4705] <= 8187;
      adc_rom[4706] <= 8188;
      adc_rom[4707] <= 8189;
      adc_rom[4708] <= 8186;
      adc_rom[4709] <= 8188;
      adc_rom[4710] <= 8185;
      adc_rom[4711] <= 8187;
      adc_rom[4712] <= 8186;
      adc_rom[4713] <= 8185;
      adc_rom[4714] <= 8187;
      adc_rom[4715] <= 8187;
      adc_rom[4716] <= 8189;
      adc_rom[4717] <= 8188;
      adc_rom[4718] <= 8185;
      adc_rom[4719] <= 8187;
      adc_rom[4720] <= 8186;
      adc_rom[4721] <= 8188;
      adc_rom[4722] <= 8187;
      adc_rom[4723] <= 8184;
      adc_rom[4724] <= 8187;
      adc_rom[4725] <= 8185;
      adc_rom[4726] <= 8187;
      adc_rom[4727] <= 8189;
      adc_rom[4728] <= 8185;
      adc_rom[4729] <= 8186;
      adc_rom[4730] <= 8186;
      adc_rom[4731] <= 8187;
      adc_rom[4732] <= 8189;
      adc_rom[4733] <= 8187;
      adc_rom[4734] <= 8187;
      adc_rom[4735] <= 8186;
      adc_rom[4736] <= 8187;
      adc_rom[4737] <= 8187;
      adc_rom[4738] <= 8185;
      adc_rom[4739] <= 8189;
      adc_rom[4740] <= 8188;
      adc_rom[4741] <= 8186;
      adc_rom[4742] <= 8187;
      adc_rom[4743] <= 8186;
      adc_rom[4744] <= 8189;
      adc_rom[4745] <= 8187;
      adc_rom[4746] <= 8187;
      adc_rom[4747] <= 8187;
      adc_rom[4748] <= 8186;
      adc_rom[4749] <= 8187;
      adc_rom[4750] <= 8185;
      adc_rom[4751] <= 8187;
      adc_rom[4752] <= 8188;
      adc_rom[4753] <= 8185;
      adc_rom[4754] <= 8188;
      adc_rom[4755] <= 8189;
      adc_rom[4756] <= 8187;
      adc_rom[4757] <= 8188;
      adc_rom[4758] <= 8187;
      adc_rom[4759] <= 8186;
      adc_rom[4760] <= 8186;
      adc_rom[4761] <= 8186;
      adc_rom[4762] <= 8187;
      adc_rom[4763] <= 8187;
      adc_rom[4764] <= 8188;
      adc_rom[4765] <= 8186;
      adc_rom[4766] <= 8185;
      adc_rom[4767] <= 8189;
      adc_rom[4768] <= 8187;
      adc_rom[4769] <= 8188;
      adc_rom[4770] <= 8185;
      adc_rom[4771] <= 8188;
      adc_rom[4772] <= 8186;
      adc_rom[4773] <= 8186;
      adc_rom[4774] <= 8188;
      adc_rom[4775] <= 8185;
      adc_rom[4776] <= 8188;
      adc_rom[4777] <= 8188;
      adc_rom[4778] <= 8185;
      adc_rom[4779] <= 8187;
      adc_rom[4780] <= 8187;
      adc_rom[4781] <= 8187;
      adc_rom[4782] <= 8187;
      adc_rom[4783] <= 8188;
      adc_rom[4784] <= 8187;
      adc_rom[4785] <= 8186;
      adc_rom[4786] <= 8186;
      adc_rom[4787] <= 8187;
      adc_rom[4788] <= 8186;
      adc_rom[4789] <= 8185;
      adc_rom[4790] <= 8186;
      adc_rom[4791] <= 8187;
      adc_rom[4792] <= 8187;
      adc_rom[4793] <= 8187;
      adc_rom[4794] <= 8189;
      adc_rom[4795] <= 8185;
      adc_rom[4796] <= 8185;
      adc_rom[4797] <= 8186;
      adc_rom[4798] <= 8186;
      adc_rom[4799] <= 8187;
      adc_rom[4800] <= 8185;
      adc_rom[4801] <= 8187;
      adc_rom[4802] <= 8187;
      adc_rom[4803] <= 8186;
      adc_rom[4804] <= 8189;
      adc_rom[4805] <= 8187;
      adc_rom[4806] <= 8187;
      adc_rom[4807] <= 8187;
      adc_rom[4808] <= 8186;
      adc_rom[4809] <= 8186;
      adc_rom[4810] <= 8186;
      adc_rom[4811] <= 8187;
      adc_rom[4812] <= 8185;
      adc_rom[4813] <= 8185;
      adc_rom[4814] <= 8187;
      adc_rom[4815] <= 8186;
      adc_rom[4816] <= 8186;
      adc_rom[4817] <= 8186;
      adc_rom[4818] <= 8185;
      adc_rom[4819] <= 8188;
      adc_rom[4820] <= 8187;
      adc_rom[4821] <= 8187;
      adc_rom[4822] <= 8187;
      adc_rom[4823] <= 8186;
      adc_rom[4824] <= 8188;
      adc_rom[4825] <= 8186;
      adc_rom[4826] <= 8186;
      adc_rom[4827] <= 8187;
      adc_rom[4828] <= 8185;
      adc_rom[4829] <= 8189;
      adc_rom[4830] <= 8185;
      adc_rom[4831] <= 8188;
      adc_rom[4832] <= 8186;
      adc_rom[4833] <= 8184;
      adc_rom[4834] <= 8187;
      adc_rom[4835] <= 8186;
      adc_rom[4836] <= 8186;
      adc_rom[4837] <= 8187;
      adc_rom[4838] <= 8186;
      adc_rom[4839] <= 8187;
      adc_rom[4840] <= 8187;
      adc_rom[4841] <= 8187;
      adc_rom[4842] <= 8189;
      adc_rom[4843] <= 8186;
      adc_rom[4844] <= 8188;
      adc_rom[4845] <= 8188;
      adc_rom[4846] <= 8185;
      adc_rom[4847] <= 8185;
      adc_rom[4848] <= 8186;
      adc_rom[4849] <= 8186;
      adc_rom[4850] <= 8188;
      adc_rom[4851] <= 8186;
      adc_rom[4852] <= 8186;
      adc_rom[4853] <= 8185;
      adc_rom[4854] <= 8187;
      adc_rom[4855] <= 8187;
      adc_rom[4856] <= 8187;
      adc_rom[4857] <= 8186;
      adc_rom[4858] <= 8185;
      adc_rom[4859] <= 8187;
      adc_rom[4860] <= 8186;
      adc_rom[4861] <= 8187;
      adc_rom[4862] <= 8187;
      adc_rom[4863] <= 8187;
      adc_rom[4864] <= 8187;
      adc_rom[4865] <= 8187;
      adc_rom[4866] <= 8189;
      adc_rom[4867] <= 8188;
      adc_rom[4868] <= 8185;
      adc_rom[4869] <= 8187;
      adc_rom[4870] <= 8187;
      adc_rom[4871] <= 8184;
      adc_rom[4872] <= 8189;
      adc_rom[4873] <= 8185;
      adc_rom[4874] <= 8187;
      adc_rom[4875] <= 8184;
      adc_rom[4876] <= 8188;
      adc_rom[4877] <= 8188;
      adc_rom[4878] <= 8186;
      adc_rom[4879] <= 8187;
      adc_rom[4880] <= 8186;
      adc_rom[4881] <= 8187;
      adc_rom[4882] <= 8187;
      adc_rom[4883] <= 8186;
      adc_rom[4884] <= 8186;
      adc_rom[4885] <= 8185;
      adc_rom[4886] <= 8184;
      adc_rom[4887] <= 8186;
      adc_rom[4888] <= 8184;
      adc_rom[4889] <= 8187;
      adc_rom[4890] <= 8186;
      adc_rom[4891] <= 8187;
      adc_rom[4892] <= 8186;
      adc_rom[4893] <= 8185;
      adc_rom[4894] <= 8186;
      adc_rom[4895] <= 8186;
      adc_rom[4896] <= 8187;
      adc_rom[4897] <= 8190;
      adc_rom[4898] <= 8185;
      adc_rom[4899] <= 8188;
      adc_rom[4900] <= 8184;
      adc_rom[4901] <= 8187;
      adc_rom[4902] <= 8186;
      adc_rom[4903] <= 8185;
      adc_rom[4904] <= 8189;
      adc_rom[4905] <= 8186;
      adc_rom[4906] <= 8187;
      adc_rom[4907] <= 8187;
      adc_rom[4908] <= 8185;
      adc_rom[4909] <= 8189;
      adc_rom[4910] <= 8185;
      adc_rom[4911] <= 8185;
      adc_rom[4912] <= 8186;
      adc_rom[4913] <= 8185;
      adc_rom[4914] <= 8186;
      adc_rom[4915] <= 8185;
      adc_rom[4916] <= 8186;
      adc_rom[4917] <= 8188;
      adc_rom[4918] <= 8185;
      adc_rom[4919] <= 8187;
      adc_rom[4920] <= 8187;
      adc_rom[4921] <= 8185;
      adc_rom[4922] <= 8186;
      adc_rom[4923] <= 8185;
      adc_rom[4924] <= 8186;
      adc_rom[4925] <= 8187;
      adc_rom[4926] <= 8187;
      adc_rom[4927] <= 8188;
      adc_rom[4928] <= 8185;
      adc_rom[4929] <= 8187;
      adc_rom[4930] <= 8186;
      adc_rom[4931] <= 8187;
      adc_rom[4932] <= 8185;
      adc_rom[4933] <= 8186;
      adc_rom[4934] <= 8188;
      adc_rom[4935] <= 8189;
      adc_rom[4936] <= 8190;
      adc_rom[4937] <= 8187;
      adc_rom[4938] <= 8187;
      adc_rom[4939] <= 8187;
      adc_rom[4940] <= 8187;
      adc_rom[4941] <= 8186;
      adc_rom[4942] <= 8190;
      adc_rom[4943] <= 8186;
      adc_rom[4944] <= 8189;
      adc_rom[4945] <= 8188;
      adc_rom[4946] <= 8188;
      adc_rom[4947] <= 8187;
      adc_rom[4948] <= 8185;
      adc_rom[4949] <= 8188;
      adc_rom[4950] <= 8185;
      adc_rom[4951] <= 8187;
      adc_rom[4952] <= 8189;
      adc_rom[4953] <= 8186;
      adc_rom[4954] <= 8187;
      adc_rom[4955] <= 8186;
      adc_rom[4956] <= 8187;
      adc_rom[4957] <= 8187;
      adc_rom[4958] <= 8186;
      adc_rom[4959] <= 8187;
      adc_rom[4960] <= 8188;
      adc_rom[4961] <= 8189;
      adc_rom[4962] <= 8187;
      adc_rom[4963] <= 8185;
      adc_rom[4964] <= 8188;
      adc_rom[4965] <= 8188;
      adc_rom[4966] <= 8190;
      adc_rom[4967] <= 8189;
      adc_rom[4968] <= 8187;
      adc_rom[4969] <= 8189;
      adc_rom[4970] <= 8186;
      adc_rom[4971] <= 8187;
      adc_rom[4972] <= 8186;
      adc_rom[4973] <= 8186;
      adc_rom[4974] <= 8187;
      adc_rom[4975] <= 8186;
      adc_rom[4976] <= 8185;
      adc_rom[4977] <= 8187;
      adc_rom[4978] <= 8185;
      adc_rom[4979] <= 8190;
      adc_rom[4980] <= 8187;
      adc_rom[4981] <= 8185;
      adc_rom[4982] <= 8188;
      adc_rom[4983] <= 8187;
      adc_rom[4984] <= 8187;
      adc_rom[4985] <= 8186;
      adc_rom[4986] <= 8186;
      adc_rom[4987] <= 8189;
      adc_rom[4988] <= 8187;
      adc_rom[4989] <= 8187;
      adc_rom[4990] <= 8186;
      adc_rom[4991] <= 8189;
      adc_rom[4992] <= 8188;
      adc_rom[4993] <= 8186;
      adc_rom[4994] <= 8188;
      adc_rom[4995] <= 8187;
      adc_rom[4996] <= 8188;
      adc_rom[4997] <= 8187;
      adc_rom[4998] <= 8188;
      adc_rom[4999] <= 8189;
      adc_rom[5000] <= 8188;
      adc_rom[5001] <= 8187;
      adc_rom[5002] <= 8190;
      adc_rom[5003] <= 8187;
      adc_rom[5004] <= 8188;
      adc_rom[5005] <= 8187;
      adc_rom[5006] <= 8187;
      adc_rom[5007] <= 8188;
      adc_rom[5008] <= 8188;
      adc_rom[5009] <= 8187;
      adc_rom[5010] <= 8185;
      adc_rom[5011] <= 8185;
      adc_rom[5012] <= 8187;
      adc_rom[5013] <= 8186;
      adc_rom[5014] <= 8186;
      adc_rom[5015] <= 8187;
      adc_rom[5016] <= 8188;
      adc_rom[5017] <= 8190;
      adc_rom[5018] <= 8187;
      adc_rom[5019] <= 8189;
      adc_rom[5020] <= 8185;
      adc_rom[5021] <= 8189;
      adc_rom[5022] <= 8188;
      adc_rom[5023] <= 8186;
      adc_rom[5024] <= 8187;
      adc_rom[5025] <= 8186;
      adc_rom[5026] <= 8187;
      adc_rom[5027] <= 8187;
      adc_rom[5028] <= 8185;
      adc_rom[5029] <= 8189;
      adc_rom[5030] <= 8189;
      adc_rom[5031] <= 8187;
      adc_rom[5032] <= 8186;
      adc_rom[5033] <= 8187;
      adc_rom[5034] <= 8187;
      adc_rom[5035] <= 8186;
      adc_rom[5036] <= 8187;
      adc_rom[5037] <= 8190;
      adc_rom[5038] <= 8187;
      adc_rom[5039] <= 8187;
      adc_rom[5040] <= 8188;
      adc_rom[5041] <= 8186;
      adc_rom[5042] <= 8186;
      adc_rom[5043] <= 8185;
      adc_rom[5044] <= 8188;
      adc_rom[5045] <= 8186;
      adc_rom[5046] <= 8189;
      adc_rom[5047] <= 8189;
      adc_rom[5048] <= 8186;
      adc_rom[5049] <= 8186;
      adc_rom[5050] <= 8188;
      adc_rom[5051] <= 8186;
      adc_rom[5052] <= 8187;
      adc_rom[5053] <= 8184;
      adc_rom[5054] <= 8188;
      adc_rom[5055] <= 8186;
      adc_rom[5056] <= 8186;
      adc_rom[5057] <= 8187;
      adc_rom[5058] <= 8187;
      adc_rom[5059] <= 8189;
      adc_rom[5060] <= 8188;
      adc_rom[5061] <= 8187;
      adc_rom[5062] <= 8188;
      adc_rom[5063] <= 8189;
      adc_rom[5064] <= 8189;
      adc_rom[5065] <= 8187;
      adc_rom[5066] <= 8188;
      adc_rom[5067] <= 8187;
      adc_rom[5068] <= 8186;
      adc_rom[5069] <= 8187;
      adc_rom[5070] <= 8185;
      adc_rom[5071] <= 8187;
      adc_rom[5072] <= 8187;
      adc_rom[5073] <= 8186;
      adc_rom[5074] <= 8187;
      adc_rom[5075] <= 8186;
      adc_rom[5076] <= 8187;
      adc_rom[5077] <= 8187;
      adc_rom[5078] <= 8185;
      adc_rom[5079] <= 8187;
      adc_rom[5080] <= 8187;
      adc_rom[5081] <= 8187;
      adc_rom[5082] <= 8189;
      adc_rom[5083] <= 8187;
      adc_rom[5084] <= 8187;
      adc_rom[5085] <= 8187;
      adc_rom[5086] <= 8187;
      adc_rom[5087] <= 8187;
      adc_rom[5088] <= 8186;
      adc_rom[5089] <= 8187;
      adc_rom[5090] <= 8188;
      adc_rom[5091] <= 8185;
      adc_rom[5092] <= 8187;
      adc_rom[5093] <= 8185;
      adc_rom[5094] <= 8188;
      adc_rom[5095] <= 8187;
      adc_rom[5096] <= 8186;
      adc_rom[5097] <= 8186;
      adc_rom[5098] <= 8185;
      adc_rom[5099] <= 8187;
      adc_rom[5100] <= 8186;
      adc_rom[5101] <= 8188;
      adc_rom[5102] <= 8185;
      adc_rom[5103] <= 8185;
      adc_rom[5104] <= 8189;
      adc_rom[5105] <= 8186;
      adc_rom[5106] <= 8188;
      adc_rom[5107] <= 8189;
      adc_rom[5108] <= 8186;
      adc_rom[5109] <= 8187;
      adc_rom[5110] <= 8187;
      adc_rom[5111] <= 8186;
      adc_rom[5112] <= 8188;
      adc_rom[5113] <= 8186;
      adc_rom[5114] <= 8188;
      adc_rom[5115] <= 8185;
      adc_rom[5116] <= 8189;
      adc_rom[5117] <= 8187;
      adc_rom[5118] <= 8185;
      adc_rom[5119] <= 8187;
      adc_rom[5120] <= 8187;
      adc_rom[5121] <= 8187;
      adc_rom[5122] <= 8186;
      adc_rom[5123] <= 8186;
      adc_rom[5124] <= 8186;
      adc_rom[5125] <= 8185;
      adc_rom[5126] <= 8188;
      adc_rom[5127] <= 8186;
      adc_rom[5128] <= 8186;
      adc_rom[5129] <= 8189;
      adc_rom[5130] <= 8185;
      adc_rom[5131] <= 8184;
      adc_rom[5132] <= 8186;
      adc_rom[5133] <= 8186;
      adc_rom[5134] <= 8189;
      adc_rom[5135] <= 8189;
      adc_rom[5136] <= 8187;
      adc_rom[5137] <= 8187;
      adc_rom[5138] <= 8187;
      adc_rom[5139] <= 8187;
      adc_rom[5140] <= 8186;
      adc_rom[5141] <= 8185;
      adc_rom[5142] <= 8187;
      adc_rom[5143] <= 8186;
      adc_rom[5144] <= 8189;
      adc_rom[5145] <= 8186;
      adc_rom[5146] <= 8189;
      adc_rom[5147] <= 8187;
      adc_rom[5148] <= 8185;
      adc_rom[5149] <= 8187;
      adc_rom[5150] <= 8185;
      adc_rom[5151] <= 8189;
      adc_rom[5152] <= 8189;
      adc_rom[5153] <= 8186;
      adc_rom[5154] <= 8186;
      adc_rom[5155] <= 8185;
      adc_rom[5156] <= 8186;
      adc_rom[5157] <= 8188;
      adc_rom[5158] <= 8185;
      adc_rom[5159] <= 8188;
      adc_rom[5160] <= 8187;
      adc_rom[5161] <= 8186;
      adc_rom[5162] <= 8189;
      adc_rom[5163] <= 8185;
      adc_rom[5164] <= 8186;
      adc_rom[5165] <= 8187;
      adc_rom[5166] <= 8186;
      adc_rom[5167] <= 8188;
      adc_rom[5168] <= 8185;
      adc_rom[5169] <= 8186;
      adc_rom[5170] <= 8186;
      adc_rom[5171] <= 8187;
      adc_rom[5172] <= 8186;
      adc_rom[5173] <= 8186;
      adc_rom[5174] <= 8186;
      adc_rom[5175] <= 8186;
      adc_rom[5176] <= 8188;
      adc_rom[5177] <= 8187;
      adc_rom[5178] <= 8186;
      adc_rom[5179] <= 8187;
      adc_rom[5180] <= 8187;
      adc_rom[5181] <= 8184;
      adc_rom[5182] <= 8186;
      adc_rom[5183] <= 8186;
      adc_rom[5184] <= 8185;
      adc_rom[5185] <= 8185;
      adc_rom[5186] <= 8186;
      adc_rom[5187] <= 8187;
      adc_rom[5188] <= 8185;
      adc_rom[5189] <= 8187;
      adc_rom[5190] <= 8183;
      adc_rom[5191] <= 8186;
      adc_rom[5192] <= 8187;
      adc_rom[5193] <= 8186;
      adc_rom[5194] <= 8186;
      adc_rom[5195] <= 8186;
      adc_rom[5196] <= 8185;
      adc_rom[5197] <= 8186;
      adc_rom[5198] <= 8187;
      adc_rom[5199] <= 8186;
      adc_rom[5200] <= 8186;
      adc_rom[5201] <= 8187;
      adc_rom[5202] <= 8188;
      adc_rom[5203] <= 8186;
      adc_rom[5204] <= 8187;
      adc_rom[5205] <= 8185;
      adc_rom[5206] <= 8185;
      adc_rom[5207] <= 8186;
      adc_rom[5208] <= 8187;
      adc_rom[5209] <= 8187;
      adc_rom[5210] <= 8184;
      adc_rom[5211] <= 8185;
      adc_rom[5212] <= 8187;
      adc_rom[5213] <= 8187;
      adc_rom[5214] <= 8187;
      adc_rom[5215] <= 8187;
      adc_rom[5216] <= 8185;
      adc_rom[5217] <= 8185;
      adc_rom[5218] <= 8183;
      adc_rom[5219] <= 8186;
      adc_rom[5220] <= 8186;
      adc_rom[5221] <= 8186;
      adc_rom[5222] <= 8186;
      adc_rom[5223] <= 8185;
      adc_rom[5224] <= 8186;
      adc_rom[5225] <= 8186;
      adc_rom[5226] <= 8186;
      adc_rom[5227] <= 8185;
      adc_rom[5228] <= 8185;
      adc_rom[5229] <= 8187;
      adc_rom[5230] <= 8186;
      adc_rom[5231] <= 8187;
      adc_rom[5232] <= 8187;
      adc_rom[5233] <= 8185;
      adc_rom[5234] <= 8185;
      adc_rom[5235] <= 8185;
      adc_rom[5236] <= 8185;
      adc_rom[5237] <= 8188;
      adc_rom[5238] <= 8186;
      adc_rom[5239] <= 8188;
      adc_rom[5240] <= 8186;
      adc_rom[5241] <= 8183;
      adc_rom[5242] <= 8186;
      adc_rom[5243] <= 8185;
      adc_rom[5244] <= 8186;
      adc_rom[5245] <= 8186;
      adc_rom[5246] <= 8185;
      adc_rom[5247] <= 8187;
      adc_rom[5248] <= 8186;
      adc_rom[5249] <= 8187;
      adc_rom[5250] <= 8187;
      adc_rom[5251] <= 8186;
      adc_rom[5252] <= 8187;
      adc_rom[5253] <= 8186;
      adc_rom[5254] <= 8185;
      adc_rom[5255] <= 8186;
      adc_rom[5256] <= 8187;
      adc_rom[5257] <= 8188;
      adc_rom[5258] <= 8184;
      adc_rom[5259] <= 8185;
      adc_rom[5260] <= 8185;
      adc_rom[5261] <= 8186;
      adc_rom[5262] <= 8187;
      adc_rom[5263] <= 8186;
      adc_rom[5264] <= 8186;
      adc_rom[5265] <= 8186;
      adc_rom[5266] <= 8186;
      adc_rom[5267] <= 8185;
      adc_rom[5268] <= 8186;
      adc_rom[5269] <= 8187;
      adc_rom[5270] <= 8186;
      adc_rom[5271] <= 8185;
      adc_rom[5272] <= 8187;
      adc_rom[5273] <= 8185;
      adc_rom[5274] <= 8188;
      adc_rom[5275] <= 8186;
      adc_rom[5276] <= 8187;
      adc_rom[5277] <= 8187;
      adc_rom[5278] <= 8186;
      adc_rom[5279] <= 8187;
      adc_rom[5280] <= 8187;
      adc_rom[5281] <= 8185;
      adc_rom[5282] <= 8189;
      adc_rom[5283] <= 8185;
      adc_rom[5284] <= 8187;
      adc_rom[5285] <= 8186;
      adc_rom[5286] <= 8185;
      adc_rom[5287] <= 8189;
      adc_rom[5288] <= 8186;
      adc_rom[5289] <= 8186;
      adc_rom[5290] <= 8185;
      adc_rom[5291] <= 8186;
      adc_rom[5292] <= 8187;
      adc_rom[5293] <= 8185;
      adc_rom[5294] <= 8187;
      adc_rom[5295] <= 8186;
      adc_rom[5296] <= 8186;
      adc_rom[5297] <= 8186;
      adc_rom[5298] <= 8186;
      adc_rom[5299] <= 8188;
      adc_rom[5300] <= 8185;
      adc_rom[5301] <= 8186;
      adc_rom[5302] <= 8186;
      adc_rom[5303] <= 8186;
      adc_rom[5304] <= 8187;
      adc_rom[5305] <= 8185;
      adc_rom[5306] <= 8186;
      adc_rom[5307] <= 8188;
      adc_rom[5308] <= 8185;
      adc_rom[5309] <= 8187;
      adc_rom[5310] <= 8185;
      adc_rom[5311] <= 8187;
      adc_rom[5312] <= 8187;
      adc_rom[5313] <= 8183;
      adc_rom[5314] <= 8188;
      adc_rom[5315] <= 8189;
      adc_rom[5316] <= 8187;
      adc_rom[5317] <= 8186;
      adc_rom[5318] <= 8183;
      adc_rom[5319] <= 8187;
      adc_rom[5320] <= 8186;
      adc_rom[5321] <= 8186;
      adc_rom[5322] <= 8189;
      adc_rom[5323] <= 8185;
      adc_rom[5324] <= 8187;
      adc_rom[5325] <= 8187;
      adc_rom[5326] <= 8187;
      adc_rom[5327] <= 8185;
      adc_rom[5328] <= 8186;
      adc_rom[5329] <= 8187;
      adc_rom[5330] <= 8186;
      adc_rom[5331] <= 8186;
      adc_rom[5332] <= 8187;
      adc_rom[5333] <= 8186;
      adc_rom[5334] <= 8187;
      adc_rom[5335] <= 8187;
      adc_rom[5336] <= 8186;
      adc_rom[5337] <= 8188;
      adc_rom[5338] <= 8184;
      adc_rom[5339] <= 8188;
      adc_rom[5340] <= 8185;
      adc_rom[5341] <= 8187;
      adc_rom[5342] <= 8188;
      adc_rom[5343] <= 8185;
      adc_rom[5344] <= 8188;
      adc_rom[5345] <= 8185;
      adc_rom[5346] <= 8187;
      adc_rom[5347] <= 8187;
      adc_rom[5348] <= 8186;
      adc_rom[5349] <= 8190;
      adc_rom[5350] <= 8185;
      adc_rom[5351] <= 8186;
      adc_rom[5352] <= 8188;
      adc_rom[5353] <= 8186;
      adc_rom[5354] <= 8188;
      adc_rom[5355] <= 8185;
      adc_rom[5356] <= 8186;
      adc_rom[5357] <= 8186;
      adc_rom[5358] <= 8184;
      adc_rom[5359] <= 8185;
      adc_rom[5360] <= 8186;
      adc_rom[5361] <= 8188;
      adc_rom[5362] <= 8186;
      adc_rom[5363] <= 8184;
      adc_rom[5364] <= 8188;
      adc_rom[5365] <= 8187;
      adc_rom[5366] <= 8186;
      adc_rom[5367] <= 8186;
      adc_rom[5368] <= 8185;
      adc_rom[5369] <= 8188;
      adc_rom[5370] <= 8185;
      adc_rom[5371] <= 8186;
      adc_rom[5372] <= 8188;
      adc_rom[5373] <= 8186;
      adc_rom[5374] <= 8189;
      adc_rom[5375] <= 8187;
      adc_rom[5376] <= 8186;
      adc_rom[5377] <= 8187;
      adc_rom[5378] <= 8186;
      adc_rom[5379] <= 8186;
      adc_rom[5380] <= 8188;
      adc_rom[5381] <= 8185;
      adc_rom[5382] <= 8188;
      adc_rom[5383] <= 8187;
      adc_rom[5384] <= 8187;
      adc_rom[5385] <= 8185;
      adc_rom[5386] <= 8186;
      adc_rom[5387] <= 8185;
      adc_rom[5388] <= 8185;
      adc_rom[5389] <= 8188;
      adc_rom[5390] <= 8186;
      adc_rom[5391] <= 8187;
      adc_rom[5392] <= 8187;
      adc_rom[5393] <= 8184;
      adc_rom[5394] <= 8188;
      adc_rom[5395] <= 8187;
      adc_rom[5396] <= 8187;
      adc_rom[5397] <= 8186;
      adc_rom[5398] <= 8185;
      adc_rom[5399] <= 8187;
      adc_rom[5400] <= 8187;
      adc_rom[5401] <= 8187;
      adc_rom[5402] <= 8187;
      adc_rom[5403] <= 8187;
      adc_rom[5404] <= 8188;
      adc_rom[5405] <= 8187;
      adc_rom[5406] <= 8187;
      adc_rom[5407] <= 8187;
      adc_rom[5408] <= 8186;
      adc_rom[5409] <= 8188;
      adc_rom[5410] <= 8185;
      adc_rom[5411] <= 8187;
      adc_rom[5412] <= 8188;
      adc_rom[5413] <= 8186;
      adc_rom[5414] <= 8188;
      adc_rom[5415] <= 8185;
      adc_rom[5416] <= 8187;
      adc_rom[5417] <= 8187;
      adc_rom[5418] <= 8186;
      adc_rom[5419] <= 8184;
      adc_rom[5420] <= 8187;
      adc_rom[5421] <= 8186;
      adc_rom[5422] <= 8187;
      adc_rom[5423] <= 8186;
      adc_rom[5424] <= 8186;
      adc_rom[5425] <= 8188;
      adc_rom[5426] <= 8186;
      adc_rom[5427] <= 8186;
      adc_rom[5428] <= 8187;
      adc_rom[5429] <= 8185;
      adc_rom[5430] <= 8185;
      adc_rom[5431] <= 8185;
      adc_rom[5432] <= 8186;
      adc_rom[5433] <= 8185;
      adc_rom[5434] <= 8187;
      adc_rom[5435] <= 8186;
      adc_rom[5436] <= 8187;
      adc_rom[5437] <= 8186;
      adc_rom[5438] <= 8186;
      adc_rom[5439] <= 8187;
      adc_rom[5440] <= 8185;
      adc_rom[5441] <= 8187;
      adc_rom[5442] <= 8186;
      adc_rom[5443] <= 8186;
      adc_rom[5444] <= 8186;
      adc_rom[5445] <= 8185;
      adc_rom[5446] <= 8186;
      adc_rom[5447] <= 8186;
      adc_rom[5448] <= 8185;
      adc_rom[5449] <= 8187;
      adc_rom[5450] <= 8185;
      adc_rom[5451] <= 8186;
      adc_rom[5452] <= 8186;
      adc_rom[5453] <= 8185;
      adc_rom[5454] <= 8187;
      adc_rom[5455] <= 8186;
      adc_rom[5456] <= 8187;
      adc_rom[5457] <= 8187;
      adc_rom[5458] <= 8185;
      adc_rom[5459] <= 8187;
      adc_rom[5460] <= 8187;
      adc_rom[5461] <= 8186;
      adc_rom[5462] <= 8189;
      adc_rom[5463] <= 8186;
      adc_rom[5464] <= 8185;
      adc_rom[5465] <= 8186;
      adc_rom[5466] <= 8186;
      adc_rom[5467] <= 8184;
      adc_rom[5468] <= 8185;
      adc_rom[5469] <= 8187;
      adc_rom[5470] <= 8187;
      adc_rom[5471] <= 8189;
      adc_rom[5472] <= 8188;
      adc_rom[5473] <= 8186;
      adc_rom[5474] <= 8187;
      adc_rom[5475] <= 8185;
      adc_rom[5476] <= 8186;
      adc_rom[5477] <= 8185;
      adc_rom[5478] <= 8186;
      adc_rom[5479] <= 8187;
      adc_rom[5480] <= 8186;
      adc_rom[5481] <= 8187;
      adc_rom[5482] <= 8186;
      adc_rom[5483] <= 8187;
      adc_rom[5484] <= 8186;
      adc_rom[5485] <= 8187;
      adc_rom[5486] <= 8188;
      adc_rom[5487] <= 8187;
      adc_rom[5488] <= 8186;
      adc_rom[5489] <= 8187;
      adc_rom[5490] <= 8185;
      adc_rom[5491] <= 8187;
      adc_rom[5492] <= 8186;
      adc_rom[5493] <= 8186;
      adc_rom[5494] <= 8187;
      adc_rom[5495] <= 8185;
      adc_rom[5496] <= 8185;
      adc_rom[5497] <= 8186;
      adc_rom[5498] <= 8184;
      adc_rom[5499] <= 8187;
      adc_rom[5500] <= 8183;
      adc_rom[5501] <= 8186;
      adc_rom[5502] <= 8187;
      adc_rom[5503] <= 8186;
      adc_rom[5504] <= 8185;
      adc_rom[5505] <= 8186;
      adc_rom[5506] <= 8186;
      adc_rom[5507] <= 8187;
      adc_rom[5508] <= 8183;
      adc_rom[5509] <= 8185;
      adc_rom[5510] <= 8186;
      adc_rom[5511] <= 8185;
      adc_rom[5512] <= 8187;
      adc_rom[5513] <= 8185;
      adc_rom[5514] <= 8187;
      adc_rom[5515] <= 8186;
      adc_rom[5516] <= 8187;
      adc_rom[5517] <= 8185;
      adc_rom[5518] <= 8186;
      adc_rom[5519] <= 8184;
      adc_rom[5520] <= 8186;
      adc_rom[5521] <= 8188;
      adc_rom[5522] <= 8187;
      adc_rom[5523] <= 8185;
      adc_rom[5524] <= 8188;
      adc_rom[5525] <= 8187;
      adc_rom[5526] <= 8186;
      adc_rom[5527] <= 8186;
      adc_rom[5528] <= 8187;
      adc_rom[5529] <= 8187;
      adc_rom[5530] <= 8185;
      adc_rom[5531] <= 8188;
      adc_rom[5532] <= 8186;
      adc_rom[5533] <= 8187;
      adc_rom[5534] <= 8188;
      adc_rom[5535] <= 8187;
      adc_rom[5536] <= 8188;
      adc_rom[5537] <= 8188;
      adc_rom[5538] <= 8184;
      adc_rom[5539] <= 8186;
      adc_rom[5540] <= 8186;
      adc_rom[5541] <= 8187;
      adc_rom[5542] <= 8187;
      adc_rom[5543] <= 8185;
      adc_rom[5544] <= 8188;
      adc_rom[5545] <= 8186;
      adc_rom[5546] <= 8187;
      adc_rom[5547] <= 8186;
      adc_rom[5548] <= 8189;
      adc_rom[5549] <= 8185;
      adc_rom[5550] <= 8185;
      adc_rom[5551] <= 8187;
      adc_rom[5552] <= 8186;
      adc_rom[5553] <= 8189;
      adc_rom[5554] <= 8185;
      adc_rom[5555] <= 8186;
      adc_rom[5556] <= 8187;
      adc_rom[5557] <= 8185;
      adc_rom[5558] <= 8187;
      adc_rom[5559] <= 8187;
      adc_rom[5560] <= 8186;
      adc_rom[5561] <= 8185;
      adc_rom[5562] <= 8185;
      adc_rom[5563] <= 8185;
      adc_rom[5564] <= 8186;
      adc_rom[5565] <= 8186;
      adc_rom[5566] <= 8187;
      adc_rom[5567] <= 8187;
      adc_rom[5568] <= 8185;
      adc_rom[5569] <= 8187;
      adc_rom[5570] <= 8185;
      adc_rom[5571] <= 8185;
      adc_rom[5572] <= 8187;
      adc_rom[5573] <= 8185;
      adc_rom[5574] <= 8185;
      adc_rom[5575] <= 8186;
      adc_rom[5576] <= 8185;
      adc_rom[5577] <= 8188;
      adc_rom[5578] <= 8186;
      adc_rom[5579] <= 8186;
      adc_rom[5580] <= 8185;
      adc_rom[5581] <= 8185;
      adc_rom[5582] <= 8186;
      adc_rom[5583] <= 8186;
      adc_rom[5584] <= 8185;
      adc_rom[5585] <= 8185;
      adc_rom[5586] <= 8188;
      adc_rom[5587] <= 8188;
      adc_rom[5588] <= 8185;
      adc_rom[5589] <= 8186;
      adc_rom[5590] <= 8185;
      adc_rom[5591] <= 8186;
      adc_rom[5592] <= 8186;
      adc_rom[5593] <= 8185;
      adc_rom[5594] <= 8186;
      adc_rom[5595] <= 8185;
      adc_rom[5596] <= 8187;
      adc_rom[5597] <= 8186;
      adc_rom[5598] <= 8185;
      adc_rom[5599] <= 8187;
      adc_rom[5600] <= 8186;
      adc_rom[5601] <= 8187;
      adc_rom[5602] <= 8187;
      adc_rom[5603] <= 8186;
      adc_rom[5604] <= 8187;
      adc_rom[5605] <= 8185;
      adc_rom[5606] <= 8186;
      adc_rom[5607] <= 8187;
      adc_rom[5608] <= 8185;
      adc_rom[5609] <= 8188;
      adc_rom[5610] <= 8183;
      adc_rom[5611] <= 8188;
      adc_rom[5612] <= 8187;
      adc_rom[5613] <= 8184;
      adc_rom[5614] <= 8186;
      adc_rom[5615] <= 8185;
      adc_rom[5616] <= 8186;
      adc_rom[5617] <= 8186;
      adc_rom[5618] <= 8186;
      adc_rom[5619] <= 8187;
      adc_rom[5620] <= 8186;
      adc_rom[5621] <= 8189;
      adc_rom[5622] <= 8186;
      adc_rom[5623] <= 8186;
      adc_rom[5624] <= 8187;
      adc_rom[5625] <= 8187;
      adc_rom[5626] <= 8186;
      adc_rom[5627] <= 8186;
      adc_rom[5628] <= 8186;
      adc_rom[5629] <= 8188;
      adc_rom[5630] <= 8185;
      adc_rom[5631] <= 8185;
      adc_rom[5632] <= 8186;
      adc_rom[5633] <= 8184;
      adc_rom[5634] <= 8186;
      adc_rom[5635] <= 8187;
      adc_rom[5636] <= 8188;
      adc_rom[5637] <= 8186;
      adc_rom[5638] <= 8185;
      adc_rom[5639] <= 8189;
      adc_rom[5640] <= 8185;
      adc_rom[5641] <= 8187;
      adc_rom[5642] <= 8188;
      adc_rom[5643] <= 8184;
      adc_rom[5644] <= 8187;
      adc_rom[5645] <= 8187;
      adc_rom[5646] <= 8186;
      adc_rom[5647] <= 8186;
      adc_rom[5648] <= 8186;
      adc_rom[5649] <= 8188;
      adc_rom[5650] <= 8188;
      adc_rom[5651] <= 8187;
      adc_rom[5652] <= 8187;
      adc_rom[5653] <= 8185;
      adc_rom[5654] <= 8186;
      adc_rom[5655] <= 8187;
      adc_rom[5656] <= 8186;
      adc_rom[5657] <= 8186;
      adc_rom[5658] <= 8187;
      adc_rom[5659] <= 8187;
      adc_rom[5660] <= 8186;
      adc_rom[5661] <= 8187;
      adc_rom[5662] <= 8185;
      adc_rom[5663] <= 8185;
      adc_rom[5664] <= 8188;
      adc_rom[5665] <= 8184;
      adc_rom[5666] <= 8189;
      adc_rom[5667] <= 8187;
      adc_rom[5668] <= 8183;
      adc_rom[5669] <= 8187;
      adc_rom[5670] <= 8185;
      adc_rom[5671] <= 8186;
      adc_rom[5672] <= 8187;
      adc_rom[5673] <= 8187;
      adc_rom[5674] <= 8189;
      adc_rom[5675] <= 8186;
      adc_rom[5676] <= 8185;
      adc_rom[5677] <= 8186;
      adc_rom[5678] <= 8187;
      adc_rom[5679] <= 8188;
      adc_rom[5680] <= 8186;
      adc_rom[5681] <= 8190;
      adc_rom[5682] <= 8188;
      adc_rom[5683] <= 8183;
      adc_rom[5684] <= 8186;
      adc_rom[5685] <= 8187;
      adc_rom[5686] <= 8188;
      adc_rom[5687] <= 8187;
      adc_rom[5688] <= 8185;
      adc_rom[5689] <= 8187;
      adc_rom[5690] <= 8186;
      adc_rom[5691] <= 8186;
      adc_rom[5692] <= 8185;
      adc_rom[5693] <= 8186;
      adc_rom[5694] <= 8188;
      adc_rom[5695] <= 8185;
      adc_rom[5696] <= 8187;
      adc_rom[5697] <= 8188;
      adc_rom[5698] <= 8187;
      adc_rom[5699] <= 8188;
      adc_rom[5700] <= 8186;
      adc_rom[5701] <= 8189;
      adc_rom[5702] <= 8187;
      adc_rom[5703] <= 8185;
      adc_rom[5704] <= 8186;
      adc_rom[5705] <= 8186;
      adc_rom[5706] <= 8187;
      adc_rom[5707] <= 8188;
      adc_rom[5708] <= 8186;
      adc_rom[5709] <= 8186;
      adc_rom[5710] <= 8187;
      adc_rom[5711] <= 8189;
      adc_rom[5712] <= 8187;
      adc_rom[5713] <= 8186;
      adc_rom[5714] <= 8189;
      adc_rom[5715] <= 8184;
      adc_rom[5716] <= 8186;
      adc_rom[5717] <= 8187;
      adc_rom[5718] <= 8184;
      adc_rom[5719] <= 8186;
      adc_rom[5720] <= 8185;
      adc_rom[5721] <= 8186;
      adc_rom[5722] <= 8185;
      adc_rom[5723] <= 8185;
      adc_rom[5724] <= 8187;
      adc_rom[5725] <= 8186;
      adc_rom[5726] <= 8187;
      adc_rom[5727] <= 8187;
      adc_rom[5728] <= 8185;
      adc_rom[5729] <= 8187;
      adc_rom[5730] <= 8185;
      adc_rom[5731] <= 8187;
      adc_rom[5732] <= 8189;
      adc_rom[5733] <= 8185;
      adc_rom[5734] <= 8188;
      adc_rom[5735] <= 8187;
      adc_rom[5736] <= 8185;
      adc_rom[5737] <= 8187;
      adc_rom[5738] <= 8186;
      adc_rom[5739] <= 8188;
      adc_rom[5740] <= 8186;
      adc_rom[5741] <= 8187;
      adc_rom[5742] <= 8187;
      adc_rom[5743] <= 8187;
      adc_rom[5744] <= 8186;
      adc_rom[5745] <= 8185;
      adc_rom[5746] <= 8187;
      adc_rom[5747] <= 8189;
      adc_rom[5748] <= 8186;
      adc_rom[5749] <= 8188;
      adc_rom[5750] <= 8187;
      adc_rom[5751] <= 8189;
      adc_rom[5752] <= 8187;
      adc_rom[5753] <= 8185;
      adc_rom[5754] <= 8187;
      adc_rom[5755] <= 8189;
      adc_rom[5756] <= 8186;
      adc_rom[5757] <= 8189;
      adc_rom[5758] <= 8188;
      adc_rom[5759] <= 8189;
      adc_rom[5760] <= 8186;
      adc_rom[5761] <= 8186;
      adc_rom[5762] <= 8188;
      adc_rom[5763] <= 8188;
      adc_rom[5764] <= 8187;
      adc_rom[5765] <= 8186;
      adc_rom[5766] <= 8187;
      adc_rom[5767] <= 8188;
      adc_rom[5768] <= 8186;
      adc_rom[5769] <= 8189;
      adc_rom[5770] <= 8187;
      adc_rom[5771] <= 8187;
      adc_rom[5772] <= 8189;
      adc_rom[5773] <= 8186;
      adc_rom[5774] <= 8188;
      adc_rom[5775] <= 8185;
      adc_rom[5776] <= 8185;
      adc_rom[5777] <= 8186;
      adc_rom[5778] <= 8187;
      adc_rom[5779] <= 8187;
      adc_rom[5780] <= 8185;
      adc_rom[5781] <= 8188;
      adc_rom[5782] <= 8187;
      adc_rom[5783] <= 8187;
      adc_rom[5784] <= 8187;
      adc_rom[5785] <= 8185;
      adc_rom[5786] <= 8188;
      adc_rom[5787] <= 8185;
      adc_rom[5788] <= 8185;
      adc_rom[5789] <= 8188;
      adc_rom[5790] <= 8188;
      adc_rom[5791] <= 8189;
      adc_rom[5792] <= 8187;
      adc_rom[5793] <= 8187;
      adc_rom[5794] <= 8186;
      adc_rom[5795] <= 8189;
      adc_rom[5796] <= 8187;
      adc_rom[5797] <= 8186;
      adc_rom[5798] <= 8185;
      adc_rom[5799] <= 8189;
      adc_rom[5800] <= 8186;
      adc_rom[5801] <= 8187;
      adc_rom[5802] <= 8186;
      adc_rom[5803] <= 8187;
      adc_rom[5804] <= 8186;
      adc_rom[5805] <= 8186;
      adc_rom[5806] <= 8187;
      adc_rom[5807] <= 8187;
      adc_rom[5808] <= 8185;
      adc_rom[5809] <= 8187;
      adc_rom[5810] <= 8184;
      adc_rom[5811] <= 8187;
      adc_rom[5812] <= 8188;
      adc_rom[5813] <= 8186;
      adc_rom[5814] <= 8186;
      adc_rom[5815] <= 8187;
      adc_rom[5816] <= 8187;
      adc_rom[5817] <= 8187;
      adc_rom[5818] <= 8186;
      adc_rom[5819] <= 8189;
      adc_rom[5820] <= 8186;
      adc_rom[5821] <= 8187;
      adc_rom[5822] <= 8186;
      adc_rom[5823] <= 8185;
      adc_rom[5824] <= 8189;
      adc_rom[5825] <= 8186;
      adc_rom[5826] <= 8186;
      adc_rom[5827] <= 8188;
      adc_rom[5828] <= 8186;
      adc_rom[5829] <= 8188;
      adc_rom[5830] <= 8187;
      adc_rom[5831] <= 8189;
      adc_rom[5832] <= 8188;
      adc_rom[5833] <= 8185;
      adc_rom[5834] <= 8189;
      adc_rom[5835] <= 8186;
      adc_rom[5836] <= 8186;
      adc_rom[5837] <= 8186;
      adc_rom[5838] <= 8186;
      adc_rom[5839] <= 8187;
      adc_rom[5840] <= 8188;
      adc_rom[5841] <= 8187;
      adc_rom[5842] <= 8187;
      adc_rom[5843] <= 8187;
      adc_rom[5844] <= 8189;
      adc_rom[5845] <= 8187;
      adc_rom[5846] <= 8188;
      adc_rom[5847] <= 8186;
      adc_rom[5848] <= 8186;
      adc_rom[5849] <= 8187;
      adc_rom[5850] <= 8187;
      adc_rom[5851] <= 8185;
      adc_rom[5852] <= 8189;
      adc_rom[5853] <= 8188;
      adc_rom[5854] <= 8187;
      adc_rom[5855] <= 8187;
      adc_rom[5856] <= 8187;
      adc_rom[5857] <= 8186;
      adc_rom[5858] <= 8184;
      adc_rom[5859] <= 8187;
      adc_rom[5860] <= 8185;
      adc_rom[5861] <= 8187;
      adc_rom[5862] <= 8185;
      adc_rom[5863] <= 8187;
      adc_rom[5864] <= 8187;
      adc_rom[5865] <= 8188;
      adc_rom[5866] <= 8185;
      adc_rom[5867] <= 8187;
      adc_rom[5868] <= 8187;
      adc_rom[5869] <= 8187;
      adc_rom[5870] <= 8187;
      adc_rom[5871] <= 8186;
      adc_rom[5872] <= 8187;
      adc_rom[5873] <= 8187;
      adc_rom[5874] <= 8187;
      adc_rom[5875] <= 8185;
      adc_rom[5876] <= 8185;
      adc_rom[5877] <= 8189;
      adc_rom[5878] <= 8186;
      adc_rom[5879] <= 8185;
      adc_rom[5880] <= 8187;
      adc_rom[5881] <= 8187;
      adc_rom[5882] <= 8186;
      adc_rom[5883] <= 8186;
      adc_rom[5884] <= 8188;
      adc_rom[5885] <= 8187;
      adc_rom[5886] <= 8187;
      adc_rom[5887] <= 8187;
      adc_rom[5888] <= 8185;
      adc_rom[5889] <= 8189;
      adc_rom[5890] <= 8184;
      adc_rom[5891] <= 8189;
      adc_rom[5892] <= 8188;
      adc_rom[5893] <= 8187;
      adc_rom[5894] <= 8187;
      adc_rom[5895] <= 8187;
      adc_rom[5896] <= 8187;
      adc_rom[5897] <= 8187;
      adc_rom[5898] <= 8188;
      adc_rom[5899] <= 8187;
      adc_rom[5900] <= 8186;
      adc_rom[5901] <= 8186;
      adc_rom[5902] <= 8186;
      adc_rom[5903] <= 8185;
      adc_rom[5904] <= 8187;
      adc_rom[5905] <= 8185;
      adc_rom[5906] <= 8188;
      adc_rom[5907] <= 8187;
      adc_rom[5908] <= 8185;
      adc_rom[5909] <= 8187;
      adc_rom[5910] <= 8187;
      adc_rom[5911] <= 8188;
      adc_rom[5912] <= 8187;
      adc_rom[5913] <= 8187;
      adc_rom[5914] <= 8187;
      adc_rom[5915] <= 8186;
      adc_rom[5916] <= 8186;
      adc_rom[5917] <= 8187;
      adc_rom[5918] <= 8186;
      adc_rom[5919] <= 8186;
      adc_rom[5920] <= 8185;
      adc_rom[5921] <= 8189;
      adc_rom[5922] <= 8188;
      adc_rom[5923] <= 8187;
      adc_rom[5924] <= 8187;
      adc_rom[5925] <= 8187;
      adc_rom[5926] <= 8189;
      adc_rom[5927] <= 8187;
      adc_rom[5928] <= 8183;
      adc_rom[5929] <= 8186;
      adc_rom[5930] <= 8187;
      adc_rom[5931] <= 8189;
      adc_rom[5932] <= 8186;
      adc_rom[5933] <= 8184;
      adc_rom[5934] <= 8188;
      adc_rom[5935] <= 8186;
      adc_rom[5936] <= 8188;
      adc_rom[5937] <= 8188;
      adc_rom[5938] <= 8187;
      adc_rom[5939] <= 8187;
      adc_rom[5940] <= 8187;
      adc_rom[5941] <= 8186;
      adc_rom[5942] <= 8189;
      adc_rom[5943] <= 8185;
      adc_rom[5944] <= 8186;
      adc_rom[5945] <= 8186;
      adc_rom[5946] <= 8187;
      adc_rom[5947] <= 8187;
      adc_rom[5948] <= 8185;
      adc_rom[5949] <= 8187;
      adc_rom[5950] <= 8185;
      adc_rom[5951] <= 8187;
      adc_rom[5952] <= 8189;
      adc_rom[5953] <= 8186;
      adc_rom[5954] <= 8188;
      adc_rom[5955] <= 8187;
      adc_rom[5956] <= 8185;
      adc_rom[5957] <= 8186;
      adc_rom[5958] <= 8185;
      adc_rom[5959] <= 8187;
      adc_rom[5960] <= 8185;
      adc_rom[5961] <= 8186;
      adc_rom[5962] <= 8187;
      adc_rom[5963] <= 8186;
      adc_rom[5964] <= 8186;
      adc_rom[5965] <= 8186;
      adc_rom[5966] <= 8185;
      adc_rom[5967] <= 8187;
      adc_rom[5968] <= 8185;
      adc_rom[5969] <= 8187;
      adc_rom[5970] <= 8186;
      adc_rom[5971] <= 8188;
      adc_rom[5972] <= 8187;
      adc_rom[5973] <= 8185;
      adc_rom[5974] <= 8190;
      adc_rom[5975] <= 8187;
      adc_rom[5976] <= 8185;
      adc_rom[5977] <= 8189;
      adc_rom[5978] <= 8186;
      adc_rom[5979] <= 8187;
      adc_rom[5980] <= 8185;
      adc_rom[5981] <= 8188;
      adc_rom[5982] <= 8186;
      adc_rom[5983] <= 8185;
      adc_rom[5984] <= 8186;
      adc_rom[5985] <= 8186;
      adc_rom[5986] <= 8186;
      adc_rom[5987] <= 8187;
      adc_rom[5988] <= 8185;
      adc_rom[5989] <= 8186;
      adc_rom[5990] <= 8184;
      adc_rom[5991] <= 8187;
      adc_rom[5992] <= 8186;
      adc_rom[5993] <= 8187;
      adc_rom[5994] <= 8187;
      adc_rom[5995] <= 8187;
      adc_rom[5996] <= 8187;
      adc_rom[5997] <= 8188;
      adc_rom[5998] <= 8186;
      adc_rom[5999] <= 8188;
      adc_rom[6000] <= 8186;
      adc_rom[6001] <= 8186;
      adc_rom[6002] <= 8186;
      adc_rom[6003] <= 8185;
      adc_rom[6004] <= 8188;
      adc_rom[6005] <= 8186;
      adc_rom[6006] <= 8187;
      adc_rom[6007] <= 8187;
      adc_rom[6008] <= 8186;
      adc_rom[6009] <= 8186;
      adc_rom[6010] <= 8187;
      adc_rom[6011] <= 8186;
      adc_rom[6012] <= 8189;
      adc_rom[6013] <= 8186;
      adc_rom[6014] <= 8185;
      adc_rom[6015] <= 8185;
      adc_rom[6016] <= 8186;
      adc_rom[6017] <= 8187;
      adc_rom[6018] <= 8184;
      adc_rom[6019] <= 8187;
      adc_rom[6020] <= 8186;
      adc_rom[6021] <= 8187;
      adc_rom[6022] <= 8187;
      adc_rom[6023] <= 8184;
      adc_rom[6024] <= 8187;
      adc_rom[6025] <= 8187;
      adc_rom[6026] <= 8185;
      adc_rom[6027] <= 8187;
      adc_rom[6028] <= 8185;
      adc_rom[6029] <= 8189;
      adc_rom[6030] <= 8187;
      adc_rom[6031] <= 8188;
      adc_rom[6032] <= 8185;
      adc_rom[6033] <= 8185;
      adc_rom[6034] <= 8189;
      adc_rom[6035] <= 8186;
      adc_rom[6036] <= 8187;
      adc_rom[6037] <= 8188;
      adc_rom[6038] <= 8186;
      adc_rom[6039] <= 8188;
      adc_rom[6040] <= 8187;
      adc_rom[6041] <= 8188;
      adc_rom[6042] <= 8187;
      adc_rom[6043] <= 8185;
      adc_rom[6044] <= 8187;
      adc_rom[6045] <= 8187;
      adc_rom[6046] <= 8189;
      adc_rom[6047] <= 8189;
      adc_rom[6048] <= 8187;
      adc_rom[6049] <= 8186;
      adc_rom[6050] <= 8187;
      adc_rom[6051] <= 8187;
      adc_rom[6052] <= 8185;
      adc_rom[6053] <= 8185;
      adc_rom[6054] <= 8186;
      adc_rom[6055] <= 8186;
      adc_rom[6056] <= 8189;
      adc_rom[6057] <= 8188;
      adc_rom[6058] <= 8184;
      adc_rom[6059] <= 8187;
      adc_rom[6060] <= 8188;
      adc_rom[6061] <= 8189;
      adc_rom[6062] <= 8185;
      adc_rom[6063] <= 8185;
      adc_rom[6064] <= 8186;
      adc_rom[6065] <= 8185;
      adc_rom[6066] <= 8185;
      adc_rom[6067] <= 8186;
      adc_rom[6068] <= 8185;
      adc_rom[6069] <= 8189;
      adc_rom[6070] <= 8186;
      adc_rom[6071] <= 8189;
      adc_rom[6072] <= 8187;
      adc_rom[6073] <= 8185;
      adc_rom[6074] <= 8185;
      adc_rom[6075] <= 8187;
      adc_rom[6076] <= 8187;
      adc_rom[6077] <= 8186;
      adc_rom[6078] <= 8186;
      adc_rom[6079] <= 8187;
      adc_rom[6080] <= 8185;
      adc_rom[6081] <= 8185;
      adc_rom[6082] <= 8187;
      adc_rom[6083] <= 8185;
      adc_rom[6084] <= 8187;
      adc_rom[6085] <= 8187;
      adc_rom[6086] <= 8186;
      adc_rom[6087] <= 8186;
      adc_rom[6088] <= 8186;
      adc_rom[6089] <= 8189;
      adc_rom[6090] <= 8186;
      adc_rom[6091] <= 8187;
      adc_rom[6092] <= 8188;
      adc_rom[6093] <= 8185;
      adc_rom[6094] <= 8188;
      adc_rom[6095] <= 8186;
      adc_rom[6096] <= 8186;
      adc_rom[6097] <= 8186;
      adc_rom[6098] <= 8184;
      adc_rom[6099] <= 8187;
      adc_rom[6100] <= 8186;
      adc_rom[6101] <= 8186;
      adc_rom[6102] <= 8186;
      adc_rom[6103] <= 8184;
      adc_rom[6104] <= 8188;
      adc_rom[6105] <= 8185;
      adc_rom[6106] <= 8187;
      adc_rom[6107] <= 8187;
      adc_rom[6108] <= 8187;
      adc_rom[6109] <= 8188;
      adc_rom[6110] <= 8186;
      adc_rom[6111] <= 8187;
      adc_rom[6112] <= 8188;
      adc_rom[6113] <= 8185;
      adc_rom[6114] <= 8186;
      adc_rom[6115] <= 8186;
      adc_rom[6116] <= 8189;
      adc_rom[6117] <= 8188;
      adc_rom[6118] <= 8186;
      adc_rom[6119] <= 8187;
      adc_rom[6120] <= 8186;
      adc_rom[6121] <= 8186;
      adc_rom[6122] <= 8187;
      adc_rom[6123] <= 8185;
      adc_rom[6124] <= 8190;
      adc_rom[6125] <= 8187;
      adc_rom[6126] <= 8187;
      adc_rom[6127] <= 8189;
      adc_rom[6128] <= 8187;
      adc_rom[6129] <= 8187;
      adc_rom[6130] <= 8187;
      adc_rom[6131] <= 8188;
      adc_rom[6132] <= 8187;
      adc_rom[6133] <= 8185;
      adc_rom[6134] <= 8187;
      adc_rom[6135] <= 8188;
      adc_rom[6136] <= 8186;
      adc_rom[6137] <= 8189;
      adc_rom[6138] <= 8187;
      adc_rom[6139] <= 8188;
      adc_rom[6140] <= 8187;
      adc_rom[6141] <= 8187;
      adc_rom[6142] <= 8186;
      adc_rom[6143] <= 8186;
      adc_rom[6144] <= 8187;
      adc_rom[6145] <= 8187;
      adc_rom[6146] <= 8188;
      adc_rom[6147] <= 8187;
      adc_rom[6148] <= 8187;
      adc_rom[6149] <= 8188;
      adc_rom[6150] <= 8185;
      adc_rom[6151] <= 8188;
      adc_rom[6152] <= 8187;
      adc_rom[6153] <= 8187;
      adc_rom[6154] <= 8188;
      adc_rom[6155] <= 8186;
      adc_rom[6156] <= 8187;
      adc_rom[6157] <= 8189;
      adc_rom[6158] <= 8185;
      adc_rom[6159] <= 8186;
      adc_rom[6160] <= 8184;
      adc_rom[6161] <= 8188;
      adc_rom[6162] <= 8189;
      adc_rom[6163] <= 8186;
      adc_rom[6164] <= 8188;
      adc_rom[6165] <= 8184;
      adc_rom[6166] <= 8186;
      adc_rom[6167] <= 8187;
      adc_rom[6168] <= 8186;
      adc_rom[6169] <= 8187;
      adc_rom[6170] <= 8186;
      adc_rom[6171] <= 8187;
      adc_rom[6172] <= 8187;
      adc_rom[6173] <= 8186;
      adc_rom[6174] <= 8186;
      adc_rom[6175] <= 8185;
      adc_rom[6176] <= 8185;
      adc_rom[6177] <= 8190;
      adc_rom[6178] <= 8186;
      adc_rom[6179] <= 8188;
      adc_rom[6180] <= 8187;
      adc_rom[6181] <= 8187;
      adc_rom[6182] <= 8188;
      adc_rom[6183] <= 8188;
      adc_rom[6184] <= 8189;
      adc_rom[6185] <= 8187;
      adc_rom[6186] <= 8188;
      adc_rom[6187] <= 8188;
      adc_rom[6188] <= 8186;
      adc_rom[6189] <= 8189;
      adc_rom[6190] <= 8186;
      adc_rom[6191] <= 8186;
      adc_rom[6192] <= 8186;
      adc_rom[6193] <= 8187;
      adc_rom[6194] <= 8186;
      adc_rom[6195] <= 8186;
      adc_rom[6196] <= 8186;
      adc_rom[6197] <= 8187;
      adc_rom[6198] <= 8185;
      adc_rom[6199] <= 8187;
      adc_rom[6200] <= 8187;
      adc_rom[6201] <= 8189;
      adc_rom[6202] <= 8187;
      adc_rom[6203] <= 8186;
      adc_rom[6204] <= 8186;
      adc_rom[6205] <= 8185;
      adc_rom[6206] <= 8185;
      adc_rom[6207] <= 8187;
      adc_rom[6208] <= 8186;
      adc_rom[6209] <= 8187;
      adc_rom[6210] <= 8186;
      adc_rom[6211] <= 8186;
      adc_rom[6212] <= 8187;
      adc_rom[6213] <= 8186;
      adc_rom[6214] <= 8187;
      adc_rom[6215] <= 8186;
      adc_rom[6216] <= 8185;
      adc_rom[6217] <= 8186;
      adc_rom[6218] <= 8185;
      adc_rom[6219] <= 8188;
      adc_rom[6220] <= 8187;
      adc_rom[6221] <= 8186;
      adc_rom[6222] <= 8184;
      adc_rom[6223] <= 8185;
      adc_rom[6224] <= 8185;
      adc_rom[6225] <= 8186;
      adc_rom[6226] <= 8186;
      adc_rom[6227] <= 8188;
      adc_rom[6228] <= 8184;
      adc_rom[6229] <= 8187;
      adc_rom[6230] <= 8188;
      adc_rom[6231] <= 8188;
      adc_rom[6232] <= 8187;
      adc_rom[6233] <= 8185;
      adc_rom[6234] <= 8188;
      adc_rom[6235] <= 8185;
      adc_rom[6236] <= 8185;
      adc_rom[6237] <= 8187;
      adc_rom[6238] <= 8186;
      adc_rom[6239] <= 8189;
      adc_rom[6240] <= 8187;
      adc_rom[6241] <= 8187;
      adc_rom[6242] <= 8187;
      adc_rom[6243] <= 8187;
      adc_rom[6244] <= 8189;
      adc_rom[6245] <= 8185;
      adc_rom[6246] <= 8187;
      adc_rom[6247] <= 8186;
      adc_rom[6248] <= 8185;
      adc_rom[6249] <= 8189;
      adc_rom[6250] <= 8184;
      adc_rom[6251] <= 8187;
      adc_rom[6252] <= 8186;
      adc_rom[6253] <= 8186;
      adc_rom[6254] <= 8186;
      adc_rom[6255] <= 8187;
      adc_rom[6256] <= 8187;
      adc_rom[6257] <= 8188;
      adc_rom[6258] <= 8184;
      adc_rom[6259] <= 8187;
      adc_rom[6260] <= 8186;
      adc_rom[6261] <= 8185;
      adc_rom[6262] <= 8184;
      adc_rom[6263] <= 8186;
      adc_rom[6264] <= 8187;
      adc_rom[6265] <= 8188;
      adc_rom[6266] <= 8186;
      adc_rom[6267] <= 8185;
      adc_rom[6268] <= 8187;
      adc_rom[6269] <= 8188;
      adc_rom[6270] <= 8185;
      adc_rom[6271] <= 8185;
      adc_rom[6272] <= 8187;
      adc_rom[6273] <= 8185;
      adc_rom[6274] <= 8187;
      adc_rom[6275] <= 8187;
      adc_rom[6276] <= 8186;
      adc_rom[6277] <= 8186;
      adc_rom[6278] <= 8184;
      adc_rom[6279] <= 8188;
      adc_rom[6280] <= 8186;
      adc_rom[6281] <= 8187;
      adc_rom[6282] <= 8186;
      adc_rom[6283] <= 8186;
      adc_rom[6284] <= 8187;
      adc_rom[6285] <= 8186;
      adc_rom[6286] <= 8188;
      adc_rom[6287] <= 8186;
      adc_rom[6288] <= 8186;
      adc_rom[6289] <= 8187;
      adc_rom[6290] <= 8186;
      adc_rom[6291] <= 8186;
      adc_rom[6292] <= 8187;
      adc_rom[6293] <= 8186;
      adc_rom[6294] <= 8186;
      adc_rom[6295] <= 8185;
      adc_rom[6296] <= 8185;
      adc_rom[6297] <= 8188;
      adc_rom[6298] <= 8188;
      adc_rom[6299] <= 8187;
      adc_rom[6300] <= 8185;
      adc_rom[6301] <= 8186;
      adc_rom[6302] <= 8185;
      adc_rom[6303] <= 8185;
      adc_rom[6304] <= 8187;
      adc_rom[6305] <= 8184;
      adc_rom[6306] <= 8187;
      adc_rom[6307] <= 8189;
      adc_rom[6308] <= 8184;
      adc_rom[6309] <= 8187;
      adc_rom[6310] <= 8185;
      adc_rom[6311] <= 8187;
      adc_rom[6312] <= 8190;
      adc_rom[6313] <= 8186;
      adc_rom[6314] <= 8187;
      adc_rom[6315] <= 8186;
      adc_rom[6316] <= 8186;
      adc_rom[6317] <= 8188;
      adc_rom[6318] <= 8187;
      adc_rom[6319] <= 8188;
      adc_rom[6320] <= 8187;
      adc_rom[6321] <= 8186;
      adc_rom[6322] <= 8187;
      adc_rom[6323] <= 8185;
      adc_rom[6324] <= 8188;
      adc_rom[6325] <= 8187;
      adc_rom[6326] <= 8188;
      adc_rom[6327] <= 8188;
      adc_rom[6328] <= 8186;
      adc_rom[6329] <= 8187;
      adc_rom[6330] <= 8186;
      adc_rom[6331] <= 8189;
      adc_rom[6332] <= 8187;
      adc_rom[6333] <= 8187;
      adc_rom[6334] <= 8187;
      adc_rom[6335] <= 8185;
      adc_rom[6336] <= 8187;
      adc_rom[6337] <= 8187;
      adc_rom[6338] <= 8185;
      adc_rom[6339] <= 8187;
      adc_rom[6340] <= 8187;
      adc_rom[6341] <= 8189;
      adc_rom[6342] <= 8188;
      adc_rom[6343] <= 8185;
      adc_rom[6344] <= 8187;
      adc_rom[6345] <= 8186;
      adc_rom[6346] <= 8187;
      adc_rom[6347] <= 8188;
      adc_rom[6348] <= 8186;
      adc_rom[6349] <= 8189;
      adc_rom[6350] <= 8187;
      adc_rom[6351] <= 8188;
      adc_rom[6352] <= 8187;
      adc_rom[6353] <= 8185;
      adc_rom[6354] <= 8186;
      adc_rom[6355] <= 8185;
      adc_rom[6356] <= 8186;
      adc_rom[6357] <= 8187;
      adc_rom[6358] <= 8185;
      adc_rom[6359] <= 8187;
      adc_rom[6360] <= 8185;
      adc_rom[6361] <= 8186;
      adc_rom[6362] <= 8186;
      adc_rom[6363] <= 8189;
      adc_rom[6364] <= 8189;
      adc_rom[6365] <= 8186;
      adc_rom[6366] <= 8186;
      adc_rom[6367] <= 8187;
      adc_rom[6368] <= 8186;
      adc_rom[6369] <= 8186;
      adc_rom[6370] <= 8186;
      adc_rom[6371] <= 8187;
      adc_rom[6372] <= 8186;
      adc_rom[6373] <= 8186;
      adc_rom[6374] <= 8188;
      adc_rom[6375] <= 8187;
      adc_rom[6376] <= 8186;
      adc_rom[6377] <= 8187;
      adc_rom[6378] <= 8186;
      adc_rom[6379] <= 8188;
      adc_rom[6380] <= 8186;
      adc_rom[6381] <= 8188;
      adc_rom[6382] <= 8186;
      adc_rom[6383] <= 8186;
      adc_rom[6384] <= 8186;
      adc_rom[6385] <= 8185;
      adc_rom[6386] <= 8187;
      adc_rom[6387] <= 8187;
      adc_rom[6388] <= 8186;
      adc_rom[6389] <= 8186;
      adc_rom[6390] <= 8185;
      adc_rom[6391] <= 8187;
      adc_rom[6392] <= 8189;
      adc_rom[6393] <= 8186;
      adc_rom[6394] <= 8187;
      adc_rom[6395] <= 8188;
      adc_rom[6396] <= 8189;
      adc_rom[6397] <= 8186;
      adc_rom[6398] <= 8186;
      adc_rom[6399] <= 8186;
      adc_rom[6400] <= 8187;
      adc_rom[6401] <= 8186;
      adc_rom[6402] <= 8188;
      adc_rom[6403] <= 8186;
      adc_rom[6404] <= 8187;
      adc_rom[6405] <= 8186;
      adc_rom[6406] <= 8185;
      adc_rom[6407] <= 8188;
      adc_rom[6408] <= 8185;
      adc_rom[6409] <= 8186;
      adc_rom[6410] <= 8184;
      adc_rom[6411] <= 8187;
      adc_rom[6412] <= 8187;
      adc_rom[6413] <= 8186;
      adc_rom[6414] <= 8187;
      adc_rom[6415] <= 8188;
      adc_rom[6416] <= 8188;
      adc_rom[6417] <= 8186;
      adc_rom[6418] <= 8183;
      adc_rom[6419] <= 8187;
      adc_rom[6420] <= 8187;
      adc_rom[6421] <= 8188;
      adc_rom[6422] <= 8186;
      adc_rom[6423] <= 8189;
      adc_rom[6424] <= 8188;
      adc_rom[6425] <= 8186;
      adc_rom[6426] <= 8186;
      adc_rom[6427] <= 8188;
      adc_rom[6428] <= 8186;
      adc_rom[6429] <= 8184;
      adc_rom[6430] <= 8185;
      adc_rom[6431] <= 8186;
      adc_rom[6432] <= 8188;
      adc_rom[6433] <= 8185;
      adc_rom[6434] <= 8187;
      adc_rom[6435] <= 8187;
      adc_rom[6436] <= 8186;
      adc_rom[6437] <= 8186;
      adc_rom[6438] <= 8187;
      adc_rom[6439] <= 8185;
      adc_rom[6440] <= 8186;
      adc_rom[6441] <= 8187;
      adc_rom[6442] <= 8186;
      adc_rom[6443] <= 8186;
      adc_rom[6444] <= 8190;
      adc_rom[6445] <= 8187;
      adc_rom[6446] <= 8185;
      adc_rom[6447] <= 8188;
      adc_rom[6448] <= 8186;
      adc_rom[6449] <= 8187;
      adc_rom[6450] <= 8186;
      adc_rom[6451] <= 8185;
      adc_rom[6452] <= 8186;
      adc_rom[6453] <= 8186;
      adc_rom[6454] <= 8188;
      adc_rom[6455] <= 8186;
      adc_rom[6456] <= 8187;
      adc_rom[6457] <= 8187;
      adc_rom[6458] <= 8186;
      adc_rom[6459] <= 8186;
      adc_rom[6460] <= 8186;
      adc_rom[6461] <= 8189;
      adc_rom[6462] <= 8188;
      adc_rom[6463] <= 8184;
      adc_rom[6464] <= 8187;
      adc_rom[6465] <= 8185;
      adc_rom[6466] <= 8187;
      adc_rom[6467] <= 8186;
      adc_rom[6468] <= 8184;
      adc_rom[6469] <= 8186;
      adc_rom[6470] <= 8185;
      adc_rom[6471] <= 8188;
      adc_rom[6472] <= 8188;
      adc_rom[6473] <= 8184;
      adc_rom[6474] <= 8187;
      adc_rom[6475] <= 8185;
      adc_rom[6476] <= 8186;
      adc_rom[6477] <= 8186;
      adc_rom[6478] <= 8185;
      adc_rom[6479] <= 8187;
      adc_rom[6480] <= 8186;
      adc_rom[6481] <= 8187;
      adc_rom[6482] <= 8187;
      adc_rom[6483] <= 8187;
      adc_rom[6484] <= 8186;
      adc_rom[6485] <= 8185;
      adc_rom[6486] <= 8186;
      adc_rom[6487] <= 8187;
      adc_rom[6488] <= 8184;
      adc_rom[6489] <= 8186;
      adc_rom[6490] <= 8185;
      adc_rom[6491] <= 8186;
      adc_rom[6492] <= 8187;
      adc_rom[6493] <= 8187;
      adc_rom[6494] <= 8187;
      adc_rom[6495] <= 8188;
      adc_rom[6496] <= 8187;
      adc_rom[6497] <= 8187;
      adc_rom[6498] <= 8185;
      adc_rom[6499] <= 8187;
      adc_rom[6500] <= 8187;
      adc_rom[6501] <= 8186;
      adc_rom[6502] <= 8186;
      adc_rom[6503] <= 8185;
      adc_rom[6504] <= 8187;
      adc_rom[6505] <= 8185;
      adc_rom[6506] <= 8186;
      adc_rom[6507] <= 8185;
      adc_rom[6508] <= 8187;
      adc_rom[6509] <= 8187;
      adc_rom[6510] <= 8186;
      adc_rom[6511] <= 8185;
      adc_rom[6512] <= 8186;
      adc_rom[6513] <= 8184;
      adc_rom[6514] <= 8185;
      adc_rom[6515] <= 8186;
      adc_rom[6516] <= 8185;
      adc_rom[6517] <= 8189;
      adc_rom[6518] <= 8186;
      adc_rom[6519] <= 8190;
      adc_rom[6520] <= 8188;
      adc_rom[6521] <= 8187;
      adc_rom[6522] <= 8186;
      adc_rom[6523] <= 8186;
      adc_rom[6524] <= 8186;
      adc_rom[6525] <= 8186;
      adc_rom[6526] <= 8188;
      adc_rom[6527] <= 8187;
      adc_rom[6528] <= 8188;
      adc_rom[6529] <= 8186;
      adc_rom[6530] <= 8185;
      adc_rom[6531] <= 8185;
      adc_rom[6532] <= 8185;
      adc_rom[6533] <= 8187;
      adc_rom[6534] <= 8187;
      adc_rom[6535] <= 8184;
      adc_rom[6536] <= 8187;
      adc_rom[6537] <= 8185;
      adc_rom[6538] <= 8186;
      adc_rom[6539] <= 8189;
      adc_rom[6540] <= 8186;
      adc_rom[6541] <= 8186;
      adc_rom[6542] <= 8186;
      adc_rom[6543] <= 8186;
      adc_rom[6544] <= 8186;
      adc_rom[6545] <= 8185;
      adc_rom[6546] <= 8186;
      adc_rom[6547] <= 8185;
      adc_rom[6548] <= 8186;
      adc_rom[6549] <= 8188;
      adc_rom[6550] <= 8186;
      adc_rom[6551] <= 8185;
      adc_rom[6552] <= 8187;
      adc_rom[6553] <= 8186;
      adc_rom[6554] <= 8187;
      adc_rom[6555] <= 8186;
      adc_rom[6556] <= 8187;
      adc_rom[6557] <= 8187;
      adc_rom[6558] <= 8186;
      adc_rom[6559] <= 8187;
      adc_rom[6560] <= 8186;
      adc_rom[6561] <= 8187;
      adc_rom[6562] <= 8186;
      adc_rom[6563] <= 8186;
      adc_rom[6564] <= 8185;
      adc_rom[6565] <= 8186;
      adc_rom[6566] <= 8185;
      adc_rom[6567] <= 8185;
      adc_rom[6568] <= 8186;
      adc_rom[6569] <= 8187;
      adc_rom[6570] <= 8186;
      adc_rom[6571] <= 8187;
      adc_rom[6572] <= 8188;
      adc_rom[6573] <= 8185;
      adc_rom[6574] <= 8188;
      adc_rom[6575] <= 8186;
      adc_rom[6576] <= 8184;
      adc_rom[6577] <= 8185;
      adc_rom[6578] <= 8186;
      adc_rom[6579] <= 8187;
      adc_rom[6580] <= 8185;
      adc_rom[6581] <= 8186;
      adc_rom[6582] <= 8189;
      adc_rom[6583] <= 8186;
      adc_rom[6584] <= 8187;
      adc_rom[6585] <= 8187;
      adc_rom[6586] <= 8187;
      adc_rom[6587] <= 8188;
      adc_rom[6588] <= 8185;
      adc_rom[6589] <= 8187;
      adc_rom[6590] <= 8186;
      adc_rom[6591] <= 8187;
      adc_rom[6592] <= 8186;
      adc_rom[6593] <= 8186;
      adc_rom[6594] <= 8187;
      adc_rom[6595] <= 8185;
      adc_rom[6596] <= 8186;
      adc_rom[6597] <= 8186;
      adc_rom[6598] <= 8185;
      adc_rom[6599] <= 8187;
      adc_rom[6600] <= 8187;
      adc_rom[6601] <= 8185;
      adc_rom[6602] <= 8185;
      adc_rom[6603] <= 8183;
      adc_rom[6604] <= 8187;
      adc_rom[6605] <= 8186;
      adc_rom[6606] <= 8185;
      adc_rom[6607] <= 8185;
      adc_rom[6608] <= 8186;
      adc_rom[6609] <= 8186;
      adc_rom[6610] <= 8185;
      adc_rom[6611] <= 8185;
      adc_rom[6612] <= 8186;
      adc_rom[6613] <= 8186;
      adc_rom[6614] <= 8187;
      adc_rom[6615] <= 8186;
      adc_rom[6616] <= 8188;
      adc_rom[6617] <= 8185;
      adc_rom[6618] <= 8185;
      adc_rom[6619] <= 8188;
      adc_rom[6620] <= 8186;
      adc_rom[6621] <= 8188;
      adc_rom[6622] <= 8187;
      adc_rom[6623] <= 8187;
      adc_rom[6624] <= 8187;
      adc_rom[6625] <= 8185;
      adc_rom[6626] <= 8188;
      adc_rom[6627] <= 8187;
      adc_rom[6628] <= 8187;
      adc_rom[6629] <= 8187;
      adc_rom[6630] <= 8185;
      adc_rom[6631] <= 8185;
      adc_rom[6632] <= 8185;
      adc_rom[6633] <= 8184;
      adc_rom[6634] <= 8186;
      adc_rom[6635] <= 8185;
      adc_rom[6636] <= 8185;
      adc_rom[6637] <= 8185;
      adc_rom[6638] <= 8187;
      adc_rom[6639] <= 8186;
      adc_rom[6640] <= 8185;
      adc_rom[6641] <= 8185;
      adc_rom[6642] <= 8189;
      adc_rom[6643] <= 8186;
      adc_rom[6644] <= 8186;
      adc_rom[6645] <= 8185;
      adc_rom[6646] <= 8188;
      adc_rom[6647] <= 8186;
      adc_rom[6648] <= 8187;
      adc_rom[6649] <= 8188;
      adc_rom[6650] <= 8185;
      adc_rom[6651] <= 8187;
      adc_rom[6652] <= 8185;
      adc_rom[6653] <= 8186;
      adc_rom[6654] <= 8187;
      adc_rom[6655] <= 8185;
      adc_rom[6656] <= 8190;
      adc_rom[6657] <= 8186;
      adc_rom[6658] <= 8184;
      adc_rom[6659] <= 8184;
      adc_rom[6660] <= 8184;
      adc_rom[6661] <= 8187;
      adc_rom[6662] <= 8188;
      adc_rom[6663] <= 8186;
      adc_rom[6664] <= 8188;
      adc_rom[6665] <= 8185;
      adc_rom[6666] <= 8186;
      adc_rom[6667] <= 8187;
      adc_rom[6668] <= 8187;
      adc_rom[6669] <= 8190;
      adc_rom[6670] <= 8185;
      adc_rom[6671] <= 8187;
      adc_rom[6672] <= 8185;
      adc_rom[6673] <= 8187;
      adc_rom[6674] <= 8186;
      adc_rom[6675] <= 8185;
      adc_rom[6676] <= 8184;
      adc_rom[6677] <= 8186;
      adc_rom[6678] <= 8185;
      adc_rom[6679] <= 8188;
      adc_rom[6680] <= 8185;
      adc_rom[6681] <= 8186;
      adc_rom[6682] <= 8189;
      adc_rom[6683] <= 8186;
      adc_rom[6684] <= 8189;
      adc_rom[6685] <= 8186;
      adc_rom[6686] <= 8186;
      adc_rom[6687] <= 8187;
      adc_rom[6688] <= 8185;
      adc_rom[6689] <= 8187;
      adc_rom[6690] <= 8186;
      adc_rom[6691] <= 8185;
      adc_rom[6692] <= 8185;
      adc_rom[6693] <= 8187;
      adc_rom[6694] <= 8188;
      adc_rom[6695] <= 8187;
      adc_rom[6696] <= 8187;
      adc_rom[6697] <= 8187;
      adc_rom[6698] <= 8187;
      adc_rom[6699] <= 8187;
      adc_rom[6700] <= 8185;
      adc_rom[6701] <= 8186;
      adc_rom[6702] <= 8186;
      adc_rom[6703] <= 8188;
      adc_rom[6704] <= 8189;
      adc_rom[6705] <= 8187;
      adc_rom[6706] <= 8187;
      adc_rom[6707] <= 8185;
      adc_rom[6708] <= 8184;
      adc_rom[6709] <= 8187;
      adc_rom[6710] <= 8187;
      adc_rom[6711] <= 8185;
      adc_rom[6712] <= 8186;
      adc_rom[6713] <= 8185;
      adc_rom[6714] <= 8185;
      adc_rom[6715] <= 8186;
      adc_rom[6716] <= 8186;
      adc_rom[6717] <= 8187;
      adc_rom[6718] <= 8184;
      adc_rom[6719] <= 8187;
      adc_rom[6720] <= 8187;
      adc_rom[6721] <= 8188;
      adc_rom[6722] <= 8185;
      adc_rom[6723] <= 8185;
      adc_rom[6724] <= 8184;
      adc_rom[6725] <= 8186;
      adc_rom[6726] <= 8185;
      adc_rom[6727] <= 8187;
      adc_rom[6728] <= 8186;
      adc_rom[6729] <= 8187;
      adc_rom[6730] <= 8187;
      adc_rom[6731] <= 8187;
      adc_rom[6732] <= 8187;
      adc_rom[6733] <= 8186;
      adc_rom[6734] <= 8188;
      adc_rom[6735] <= 8186;
      adc_rom[6736] <= 8187;
      adc_rom[6737] <= 8186;
      adc_rom[6738] <= 8186;
      adc_rom[6739] <= 8186;
      adc_rom[6740] <= 8185;
      adc_rom[6741] <= 8187;
      adc_rom[6742] <= 8187;
      adc_rom[6743] <= 8187;
      adc_rom[6744] <= 8185;
      adc_rom[6745] <= 8185;
      adc_rom[6746] <= 8185;
      adc_rom[6747] <= 8188;
      adc_rom[6748] <= 8185;
      adc_rom[6749] <= 8186;
      adc_rom[6750] <= 8186;
      adc_rom[6751] <= 8187;
      adc_rom[6752] <= 8185;
      adc_rom[6753] <= 8186;
      adc_rom[6754] <= 8187;
      adc_rom[6755] <= 8184;
      adc_rom[6756] <= 8185;
      adc_rom[6757] <= 8187;
      adc_rom[6758] <= 8183;
      adc_rom[6759] <= 8187;
      adc_rom[6760] <= 8186;
      adc_rom[6761] <= 8186;
      adc_rom[6762] <= 8187;
      adc_rom[6763] <= 8183;
      adc_rom[6764] <= 8188;
      adc_rom[6765] <= 8186;
      adc_rom[6766] <= 8186;
      adc_rom[6767] <= 8187;
      adc_rom[6768] <= 8186;
      adc_rom[6769] <= 8187;
      adc_rom[6770] <= 8187;
      adc_rom[6771] <= 8187;
      adc_rom[6772] <= 8189;
      adc_rom[6773] <= 8185;
      adc_rom[6774] <= 8187;
      adc_rom[6775] <= 8186;
      adc_rom[6776] <= 8187;
      adc_rom[6777] <= 8186;
      adc_rom[6778] <= 8185;
      
   end
   
endmodule
