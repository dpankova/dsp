library verilog;
use verilog.vl_types.all;
entity IIR_avr_tst is
end IIR_avr_tst;
